magic
tech sky130A
timestamp 1716540843
<< nwell >>
rect -38 -39 59 55
<< nsubdiff >>
rect -19 18 31 31
rect -19 -8 -7 18
rect 17 -8 31 18
rect -19 -20 31 -8
<< nsubdiffcont >>
rect -7 -8 17 18
<< locali >>
rect -19 18 31 31
rect -19 -8 -7 18
rect 17 -8 31 18
rect -19 -20 31 -8
<< end >>
