magic
tech sky130A
timestamp 1717235020
<< metal3 >>
rect 0 2706 254 2745
rect 0 2589 62 2706
rect 190 2589 254 2706
rect 0 2540 254 2589
rect 0 -46 255 0
rect 0 -163 64 -46
rect 192 -163 255 -46
rect 0 -206 255 -163
<< via3 >>
rect 62 2589 190 2706
rect 64 -163 192 -46
<< metal4 >>
rect 0 2706 254 2745
rect 0 2589 62 2706
rect 190 2589 254 2706
rect 0 0 254 2589
rect 0 -46 255 0
rect 0 -163 64 -46
rect 192 -163 255 -46
rect 0 -206 255 -163
<< end >>
