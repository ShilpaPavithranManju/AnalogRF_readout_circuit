magic
tech sky130A
timestamp 1717240698
<< nmos >>
rect -100 -350 100 350
<< ndiff >>
rect -129 344 -100 350
rect -129 -344 -123 344
rect -106 -344 -100 344
rect -129 -350 -100 -344
rect 100 344 129 350
rect 100 -344 106 344
rect 123 -344 129 344
rect 100 -350 129 -344
<< ndiffc >>
rect -123 -344 -106 344
rect 106 -344 123 344
<< poly >>
rect -100 350 100 363
rect -100 -363 100 -350
<< locali >>
rect -123 344 -106 352
rect -123 -352 -106 -344
rect 106 344 123 352
rect 106 -352 123 -344
<< viali >>
rect -123 -344 -106 344
rect 106 -344 123 344
<< metal1 >>
rect -126 344 -103 350
rect -126 -344 -123 344
rect -106 -344 -103 344
rect -126 -350 -103 -344
rect 103 344 126 350
rect 103 -344 106 344
rect 123 -344 126 344
rect 103 -350 126 -344
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 7.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
