magic
tech sky130A
magscale 1 2
timestamp 1717233969
<< metal1 >>
rect 0 5903 400 6000
rect 0 5690 105 5903
rect 300 5690 400 5903
rect 0 3200 400 5690
rect 0 1800 400 2800
rect 0 316 400 1400
rect 0 103 101 316
rect 296 103 400 316
rect 0 0 400 103
<< via1 >>
rect 105 5690 300 5903
rect 101 103 296 316
<< metal2 >>
rect 0 5903 400 6000
rect 0 5690 105 5903
rect 300 5690 400 5903
rect 0 5600 400 5690
rect 0 316 400 400
rect 0 103 101 316
rect 296 103 400 316
rect 0 0 400 103
<< via2 >>
rect 105 5690 300 5903
rect 101 103 296 316
<< metal3 >>
rect 0 5903 400 6000
rect 0 5690 105 5903
rect 300 5690 400 5903
rect 0 5600 400 5690
rect 0 316 400 400
rect 0 103 101 316
rect 296 103 400 316
rect 0 0 400 103
<< via3 >>
rect 105 5690 300 5903
rect 101 103 296 316
<< metal4 >>
rect -5000 5600 -400 6000
rect 0 5903 400 6000
rect 0 5690 105 5903
rect 300 5690 400 5903
rect 0 5600 400 5690
rect -5000 -8400 -4600 5600
rect -3600 4200 8200 4600
rect -3600 -7000 -3200 4200
rect -2200 2800 6800 3200
rect -2200 -5400 -1800 2800
rect -800 1400 5400 1800
rect -800 -4000 -400 1400
rect 0 316 4000 400
rect 0 103 101 316
rect 296 103 4000 316
rect 0 0 4000 103
rect 400 -1 484 0
rect 3600 -4000 4000 0
rect -800 -4400 4000 -4000
rect 5000 -5400 5400 1400
rect -2200 -5800 5400 -5400
rect 6400 -7000 6800 2800
rect -3600 -7400 6800 -7000
rect 7798 -8400 8200 4200
rect -5000 -8800 8200 -8400
<< end >>
