magic
tech sky130A
timestamp 1717240698
<< nwell >>
rect -72 -1031 72 1031
<< pmos >>
rect -25 -1000 25 1000
<< pdiff >>
rect -54 994 -25 1000
rect -54 -994 -48 994
rect -31 -994 -25 994
rect -54 -1000 -25 -994
rect 25 994 54 1000
rect 25 -994 31 994
rect 48 -994 54 994
rect 25 -1000 54 -994
<< pdiffc >>
rect -48 -994 -31 994
rect 31 -994 48 994
<< poly >>
rect -25 1000 25 1013
rect -25 -1013 25 -1000
<< locali >>
rect -48 994 -31 1002
rect -48 -1002 -31 -994
rect 31 994 48 1002
rect 31 -1002 48 -994
<< viali >>
rect -48 -994 -31 994
rect 31 -994 48 994
<< metal1 >>
rect -51 994 -28 1000
rect -51 -994 -48 994
rect -31 -994 -28 994
rect -51 -1000 -28 -994
rect 28 994 51 1000
rect 28 -994 31 994
rect 48 -994 51 994
rect 28 -1000 51 -994
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
