magic
tech sky130A
magscale 1 2
timestamp 1717250560
<< nwell >>
rect 18 4968 90 4987
rect -2646 3608 -2313 3610
rect -3192 2745 -2313 3608
rect -3191 2742 -2313 2745
rect 179 3602 665 3603
rect 179 2738 1303 3602
rect 653 2736 1303 2738
<< psubdiff >>
rect -1046 4819 -313 4899
rect -1046 4368 -964 4819
rect -411 4368 -313 4819
rect -1046 4303 -313 4368
rect -1238 1501 -505 1581
rect -1238 1050 -1156 1501
rect -603 1050 -505 1501
rect -1238 985 -505 1050
<< nsubdiff >>
rect -3154 3386 -2648 3568
rect -3154 2931 -3061 3386
rect -2752 2931 -2648 3386
rect -3154 2788 -2648 2931
rect 690 3380 1196 3562
rect 690 2925 783 3380
rect 1092 2925 1196 3380
rect 690 2782 1196 2925
<< psubdiffcont >>
rect -964 4368 -411 4819
rect -1156 1050 -603 1501
<< nsubdiffcont >>
rect -3061 2931 -2752 3386
rect 783 2925 1092 3380
<< poly >>
rect 18 5037 90 5049
rect 18 5003 34 5037
rect 74 5003 90 5037
rect 18 4968 90 5003
rect -999 4142 -739 4169
rect -999 4026 -945 4142
rect -806 4026 -739 4142
rect -2291 3952 -2148 3957
rect -2291 3941 -1396 3952
rect -2291 3860 -2241 3941
rect -2165 3860 -1396 3941
rect -999 3882 -739 4026
rect -2291 3844 -1396 3860
rect -2255 3797 -1396 3844
rect -2255 3761 -1854 3797
rect -1797 3761 -1396 3797
rect -1469 1983 -1351 2025
rect -1595 1933 -1351 1983
rect -1928 1675 -1878 1785
rect -2227 1625 -1878 1675
rect -1773 1570 -1723 1783
rect -1595 1310 -1545 1933
rect -1469 1892 -1351 1933
rect -1603 1300 -1537 1310
rect -1603 1266 -1587 1300
rect -1553 1266 -1537 1300
rect -1603 1256 -1537 1266
<< polycont >>
rect 34 5003 74 5037
rect -945 4026 -806 4142
rect -2241 3860 -2165 3941
rect -1587 1266 -1553 1300
<< locali >>
rect -2994 5372 -2780 5413
rect -2996 5354 -2780 5372
rect -2996 5244 -2964 5354
rect -2816 5244 -2780 5354
rect -2996 3548 -2780 5244
rect 269 5324 503 5378
rect 269 5215 297 5324
rect 468 5215 503 5324
rect -1385 5040 90 5074
rect -2291 3952 -2148 3957
rect -2301 3941 -2148 3952
rect -2301 3860 -2241 3941
rect -2165 3860 -2148 3941
rect -2301 3844 -2148 3860
rect -2301 3738 -2267 3844
rect -1385 3731 -1351 5040
rect 18 5037 90 5040
rect 18 5003 34 5037
rect 74 5003 90 5037
rect 18 4987 90 5003
rect -322 4899 -257 4900
rect -1047 4819 -257 4899
rect -1047 4436 -964 4819
rect -1121 4402 -964 4436
rect -1121 3860 -1087 4402
rect -1047 4368 -964 4402
rect -411 4368 -257 4819
rect -1047 4305 -257 4368
rect -1047 4302 -258 4305
rect -1000 4142 -572 4169
rect -1000 4026 -945 4142
rect -806 4131 -572 4142
rect -806 4036 -692 4131
rect -600 4036 -572 4131
rect -806 4026 -572 4036
rect -1000 4001 -572 4026
rect -430 4107 -258 4302
rect -430 3999 -396 4107
rect -289 3999 -258 4107
rect -430 3976 -258 3999
rect -3134 3386 -2662 3548
rect -3134 2931 -3061 3386
rect -2752 2931 -2662 3386
rect -3134 2796 -2662 2931
rect -2301 2399 -2267 2535
rect -1385 2399 -1351 2535
rect -664 2452 -11 3859
rect 269 3541 503 5215
rect 710 3541 1182 3542
rect 121 3380 1182 3541
rect 121 2925 783 3380
rect 1092 2925 1182 3380
rect 121 2790 1182 2925
rect -2301 2365 -1964 2399
rect -1998 2300 -1964 2365
rect -1682 2365 -1351 2399
rect -1682 2298 -1648 2365
rect -1550 2188 -1342 2223
rect -1841 1724 -1806 1797
rect -1550 1724 -1515 2188
rect -1841 1689 -1515 1724
rect -1240 1581 -537 1734
rect -1240 1579 -503 1581
rect -1239 1501 -503 1579
rect -1587 1308 -1553 1316
rect -1587 1250 -1553 1259
rect -1239 1050 -1156 1501
rect -603 1050 -503 1501
rect -1239 984 -503 1050
rect -1239 979 -656 984
rect -1065 618 -656 979
rect -1065 462 -982 618
rect -763 462 -656 618
rect -1065 425 -656 462
<< viali >>
rect -2964 5244 -2816 5354
rect 297 5215 468 5324
rect -692 4036 -600 4131
rect -396 3999 -289 4107
rect -1594 1300 -1545 1308
rect -1594 1266 -1587 1300
rect -1587 1266 -1553 1300
rect -1553 1266 -1545 1300
rect -1594 1259 -1545 1266
rect -982 462 -763 618
<< metal1 >>
rect -3080 5354 561 5470
rect -3080 5244 -2964 5354
rect -2816 5324 561 5354
rect -2816 5244 297 5324
rect -3080 5215 297 5244
rect 468 5215 561 5324
rect -3080 5174 561 5215
rect -2557 1308 -2508 5174
rect -1909 2466 -1746 5174
rect -708 4131 -564 5174
rect -708 4036 -692 4131
rect -600 4036 -564 4131
rect -708 4001 -564 4036
rect -430 4107 -259 4151
rect -430 3999 -396 4107
rect -289 3999 -259 4107
rect -1600 1308 -1539 1320
rect -2557 1259 -1594 1308
rect -1545 1259 -1539 1308
rect -1600 1247 -1539 1259
rect -982 655 -718 661
rect -430 655 -259 3999
rect -3053 618 588 655
rect -3053 462 -982 618
rect -763 462 588 618
rect -3053 359 588 462
use sky130_fd_pr__nfet_01v8_LYFHMA  sky130_fd_pr__nfet_01v8_LYFHMA_0
timestamp 1717240698
transform -1 0 -1902 0 1 2048
box -108 -276 108 276
use sky130_fd_pr__pfet_01v8_LMLH7X  sky130_fd_pr__pfet_01v8_LMLH7X_0
timestamp 1717240698
transform 1 0 -1597 0 1 3135
box -294 -662 294 662
use sky130_fd_pr__nfet_01v8_LYFHMA  XM2
timestamp 1717240698
transform 1 0 -1744 0 1 2048
box -108 -276 108 276
use sky130_fd_pr__pfet_01v8_LMLH7X  XM3
timestamp 1717240698
transform -1 0 -2055 0 1 3135
box -294 -662 294 662
use sky130_fd_pr__pfet_01v8_A424KG  XM4
timestamp 1717240698
transform -1 0 53 0 1 2942
box -144 -2062 144 2062
use sky130_fd_pr__nfet_01v8_JAAG9L  XM5
timestamp 1717240698
transform 0 -1 -942 1 0 1977
box -258 -426 258 426
use sky130_fd_pr__nfet_01v8_DXAGR4  XM7
timestamp 1717240698
transform 1 0 -875 0 1 3157
box -258 -726 258 726
<< labels >>
rlabel space -2222 1628 -2181 1671 5 vinminus
rlabel space -1769 1579 -1728 1622 5 vinplus
rlabel locali -518 2517 -236 2647 5 vout
rlabel space -2867 418 -2779 578 5 vss
rlabel space -2625 5245 -2537 5405 5 vdd
<< end >>
