magic
tech sky130A
timestamp 1717240698
<< nwell >>
rect -147 -331 147 331
<< pmos >>
rect -100 -300 100 300
<< pdiff >>
rect -129 294 -100 300
rect -129 -294 -123 294
rect -106 -294 -100 294
rect -129 -300 -100 -294
rect 100 294 129 300
rect 100 -294 106 294
rect 123 -294 129 294
rect 100 -300 129 -294
<< pdiffc >>
rect -123 -294 -106 294
rect 106 -294 123 294
<< poly >>
rect -100 300 100 313
rect -100 -313 100 -300
<< locali >>
rect -123 294 -106 302
rect -123 -302 -106 -294
rect 106 294 123 302
rect 106 -302 123 -294
<< viali >>
rect -123 -294 -106 294
rect 106 -294 123 294
<< metal1 >>
rect -126 294 -103 300
rect -126 -294 -123 294
rect -106 -294 -103 294
rect -126 -300 -103 -294
rect 103 294 126 300
rect 103 -294 106 294
rect 123 -294 126 294
rect 103 -300 126 -294
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
