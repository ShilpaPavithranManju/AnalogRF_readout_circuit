magic
tech sky130A
magscale 1 2
timestamp 1717240620
<< nwell >>
rect -246 -2219 246 2219
<< pmos >>
rect -50 -2000 50 2000
<< pdiff >>
rect -108 1988 -50 2000
rect -108 -1988 -96 1988
rect -62 -1988 -50 1988
rect -108 -2000 -50 -1988
rect 50 1988 108 2000
rect 50 -1988 62 1988
rect 96 -1988 108 1988
rect 50 -2000 108 -1988
<< pdiffc >>
rect -96 -1988 -62 1988
rect 62 -1988 96 1988
<< nsubdiff >>
rect -210 2149 -114 2183
rect 114 2149 210 2183
rect -210 2087 -176 2149
rect 176 2087 210 2149
rect -210 -2149 -176 -2087
rect 176 -2149 210 -2087
rect -210 -2183 -114 -2149
rect 114 -2183 210 -2149
<< nsubdiffcont >>
rect -114 2149 114 2183
rect -210 -2087 -176 2087
rect 176 -2087 210 2087
rect -114 -2183 114 -2149
<< poly >>
rect -50 2081 50 2097
rect -50 2047 -34 2081
rect 34 2047 50 2081
rect -50 2000 50 2047
rect -50 -2047 50 -2000
rect -50 -2081 -34 -2047
rect 34 -2081 50 -2047
rect -50 -2097 50 -2081
<< polycont >>
rect -34 2047 34 2081
rect -34 -2081 34 -2047
<< locali >>
rect -210 2149 -114 2183
rect 114 2149 210 2183
rect -210 2087 -176 2149
rect 176 2087 210 2149
rect -50 2047 -34 2081
rect 34 2047 50 2081
rect -96 1988 -62 2004
rect -96 -2004 -62 -1988
rect 62 1988 96 2004
rect 62 -2004 96 -1988
rect -50 -2081 -34 -2047
rect 34 -2081 50 -2047
rect -210 -2149 -176 -2087
rect 176 -2149 210 -2087
rect -210 -2183 -114 -2149
rect 114 -2183 210 -2149
<< viali >>
rect -34 2047 34 2081
rect -96 -1988 -62 1988
rect 62 -1988 96 1988
rect -34 -2081 34 -2047
<< metal1 >>
rect -46 2081 46 2087
rect -46 2047 -34 2081
rect 34 2047 46 2081
rect -46 2041 46 2047
rect -102 1988 -56 2000
rect -102 -1988 -96 1988
rect -62 -1988 -56 1988
rect -102 -2000 -56 -1988
rect 56 1988 102 2000
rect 56 -1988 62 1988
rect 96 -1988 102 1988
rect 56 -2000 102 -1988
rect -46 -2047 46 -2041
rect -46 -2081 -34 -2047
rect 34 -2081 46 -2047
rect -46 -2087 46 -2081
<< properties >>
string FIXED_BBOX -193 -2166 193 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
