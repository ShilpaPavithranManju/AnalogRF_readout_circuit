magic
tech sky130A
magscale 1 2
timestamp 1717057377
<< nwell >>
rect -508 998 -330 1064
rect -138 1016 158 1064
rect -112 998 154 1016
rect -508 928 612 998
rect -508 729 508 928
rect -508 719 511 729
rect -508 707 518 719
rect -508 699 533 707
rect -508 684 518 699
rect -508 658 252 684
rect -508 626 108 658
rect -508 578 -344 626
rect -508 462 -500 578
rect -432 573 -395 578
rect -338 573 108 626
rect 488 624 518 684
rect -432 536 108 573
rect -338 494 108 536
rect -338 366 256 494
rect -122 360 256 366
<< psubdiff >>
rect -890 882 -744 921
rect -890 788 -849 882
rect -780 788 -744 882
rect -890 738 -744 788
<< nsubdiff >>
rect -455 799 -351 823
rect -455 749 -429 799
rect -376 749 -351 799
rect -455 721 -351 749
<< psubdiffcont >>
rect -849 788 -780 882
<< nsubdiffcont >>
rect -429 749 -376 799
<< poly >>
rect -236 1632 366 1662
rect -236 1433 -206 1632
rect 36 1572 106 1589
rect 36 1537 52 1572
rect 89 1567 106 1572
rect 89 1537 278 1567
rect 36 1533 278 1537
rect 36 1517 106 1533
rect 248 1483 278 1533
rect 336 1492 366 1632
rect 55 820 127 838
rect 55 785 75 820
rect 110 813 127 820
rect 336 813 366 865
rect 110 785 366 813
rect 55 776 366 785
rect 55 766 127 776
rect -61 719 5 733
rect -61 682 -45 719
rect -11 688 518 719
rect -11 682 5 688
rect -61 649 5 682
rect 182 640 212 688
rect 488 624 518 688
rect -234 -361 -204 76
rect -107 -33 -40 -16
rect -107 -67 -94 -33
rect -55 -67 -40 -33
rect -107 -85 -40 -67
rect -83 -196 -53 -85
rect 94 -196 124 0
rect 182 -57 212 8
rect 182 -68 256 -57
rect 182 -102 205 -68
rect 240 -102 256 -68
rect 182 -138 256 -102
rect 400 -196 430 26
rect -83 -226 430 -196
rect 180 -357 262 -337
rect 180 -361 206 -357
rect -234 -391 206 -361
rect 241 -361 262 -357
rect 488 -361 518 12
rect 241 -391 518 -361
rect 180 -424 262 -391
<< polycont >>
rect 52 1537 89 1572
rect 75 785 110 820
rect -45 682 -11 719
rect -94 -67 -55 -33
rect 205 -102 240 -68
rect 206 -391 241 -357
<< locali >>
rect 36 1572 106 1589
rect 36 1567 52 1572
rect -194 1537 52 1567
rect 89 1537 106 1572
rect -194 1533 106 1537
rect -194 1417 -160 1533
rect 36 1517 106 1533
rect -849 1274 -322 1308
rect -849 1272 -487 1274
rect -849 921 -775 1272
rect -433 934 -328 970
rect -890 882 -744 921
rect -890 788 -849 882
rect -780 788 -744 882
rect -433 823 -394 934
rect -890 738 -744 788
rect -455 799 -351 823
rect -455 749 -429 799
rect -376 749 -351 799
rect -194 813 -160 880
rect 55 820 127 838
rect 55 813 75 820
rect -194 785 75 813
rect 110 785 127 820
rect -194 777 127 785
rect 55 766 127 777
rect -846 232 -776 738
rect -455 721 -351 749
rect -61 722 5 733
rect -432 573 -395 721
rect -192 719 5 722
rect -192 686 -45 719
rect -192 612 -158 686
rect -61 682 -45 686
rect -11 682 5 719
rect -61 649 5 682
rect -432 536 -279 573
rect -846 222 -308 232
rect -845 198 -308 222
rect -192 -34 -157 94
rect -107 -33 -40 -16
rect -107 -34 -94 -33
rect -192 -67 -94 -34
rect -55 -67 -40 -33
rect -192 -69 -40 -67
rect -107 -85 -40 -69
rect 182 -68 256 -57
rect 182 -102 205 -68
rect 240 -102 256 -68
rect 182 -138 256 -102
rect 200 -337 235 -138
rect 180 -357 262 -337
rect 180 -391 206 -357
rect 241 -391 262 -357
rect 180 -424 262 -391
use inverter  inverter_0
timestamp 1716986487
transform 1 0 -280 0 1 -580
box -226 644 170 1266
use inverter  inverter_2
timestamp 1716986487
transform 1 0 -282 0 -1 2086
box -226 644 170 1266
use mux1_4  mux1_4_0
timestamp 1717047906
transform 1 0 0 0 1 0
box 0 0 612 1498
<< end >>
