magic
tech sky130A
magscale 1 2
timestamp 1716989908
<< viali >>
rect 3893 14025 3927 14059
rect 11069 14025 11103 14059
rect 12909 13957 12943 13991
rect 4169 13889 4203 13923
rect 10977 13889 11011 13923
rect 12725 13753 12759 13787
rect 10241 13345 10275 13379
rect 7297 13277 7331 13311
rect 7481 13277 7515 13311
rect 8125 13277 8159 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9321 13277 9355 13311
rect 9689 13277 9723 13311
rect 10517 13209 10551 13243
rect 7481 13141 7515 13175
rect 7941 13141 7975 13175
rect 9873 13141 9907 13175
rect 11989 13141 12023 13175
rect 11621 12937 11655 12971
rect 6545 12869 6579 12903
rect 6745 12869 6779 12903
rect 7021 12869 7055 12903
rect 5641 12801 5675 12835
rect 6101 12801 6135 12835
rect 7205 12801 7239 12835
rect 7481 12801 7515 12835
rect 9781 12801 9815 12835
rect 10701 12801 10735 12835
rect 11713 12801 11747 12835
rect 5733 12733 5767 12767
rect 7757 12733 7791 12767
rect 9229 12733 9263 12767
rect 9505 12733 9539 12767
rect 6377 12665 6411 12699
rect 9597 12665 9631 12699
rect 10609 12665 10643 12699
rect 5917 12597 5951 12631
rect 6561 12597 6595 12631
rect 7389 12597 7423 12631
rect 9965 12597 9999 12631
rect 7389 12393 7423 12427
rect 8585 12393 8619 12427
rect 9689 12393 9723 12427
rect 11897 12393 11931 12427
rect 7573 12325 7607 12359
rect 8401 12325 8435 12359
rect 9781 12325 9815 12359
rect 5089 12257 5123 12291
rect 8125 12257 8159 12291
rect 8033 12189 8067 12223
rect 8493 12189 8527 12223
rect 9137 12189 9171 12223
rect 9505 12189 9539 12223
rect 9965 12189 9999 12223
rect 10130 12189 10164 12223
rect 10241 12189 10275 12223
rect 10343 12199 10377 12233
rect 11989 12189 12023 12223
rect 5365 12121 5399 12155
rect 7205 12121 7239 12155
rect 7405 12121 7439 12155
rect 9321 12121 9355 12155
rect 9413 12121 9447 12155
rect 6837 12053 6871 12087
rect 11529 12053 11563 12087
rect 7021 11849 7055 11883
rect 7205 11849 7239 11883
rect 6653 11781 6687 11815
rect 6853 11781 6887 11815
rect 9781 11781 9815 11815
rect 4813 11713 4847 11747
rect 7297 11713 7331 11747
rect 9413 11713 9447 11747
rect 9505 11713 9539 11747
rect 9597 11713 9631 11747
rect 10057 11713 10091 11747
rect 10149 11713 10183 11747
rect 10425 11713 10459 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 12173 11713 12207 11747
rect 11345 11645 11379 11679
rect 11621 11645 11655 11679
rect 4629 11509 4663 11543
rect 6837 11509 6871 11543
rect 9229 11509 9263 11543
rect 9873 11509 9907 11543
rect 10333 11509 10367 11543
rect 11161 11509 11195 11543
rect 11253 11509 11287 11543
rect 11989 11509 12023 11543
rect 12265 11509 12299 11543
rect 6837 11305 6871 11339
rect 9045 11305 9079 11339
rect 11161 11305 11195 11339
rect 8125 11237 8159 11271
rect 3801 11169 3835 11203
rect 6193 11169 6227 11203
rect 7113 11169 7147 11203
rect 6101 11101 6135 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 7297 11101 7331 11135
rect 9229 11101 9263 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9607 11111 9641 11145
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 11989 11101 12023 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 4077 11033 4111 11067
rect 5825 11033 5859 11067
rect 8309 11033 8343 11067
rect 8493 11033 8527 11067
rect 11713 11033 11747 11067
rect 6469 10965 6503 10999
rect 11529 10965 11563 10999
rect 4721 10761 4755 10795
rect 6377 10761 6411 10795
rect 8033 10761 8067 10795
rect 10701 10761 10735 10795
rect 11897 10761 11931 10795
rect 6837 10693 6871 10727
rect 8401 10693 8435 10727
rect 9597 10693 9631 10727
rect 4629 10625 4663 10659
rect 5917 10625 5951 10659
rect 6101 10625 6135 10659
rect 6193 10625 6227 10659
rect 7849 10625 7883 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 8217 10625 8251 10659
rect 8493 10625 8527 10659
rect 9781 10625 9815 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 10425 10625 10459 10659
rect 10793 10625 10827 10659
rect 12725 10625 12759 10659
rect 7297 10557 7331 10591
rect 10885 10557 10919 10591
rect 13001 10557 13035 10591
rect 6469 10489 6503 10523
rect 9873 10489 9907 10523
rect 11161 10489 11195 10523
rect 11345 10489 11379 10523
rect 11529 10489 11563 10523
rect 12081 10489 12115 10523
rect 5917 10421 5951 10455
rect 8217 10421 8251 10455
rect 10333 10421 10367 10455
rect 11897 10421 11931 10455
rect 7021 10217 7055 10251
rect 9781 10217 9815 10251
rect 9965 10217 9999 10251
rect 10517 10217 10551 10251
rect 10885 10217 10919 10251
rect 12081 10217 12115 10251
rect 12357 10217 12391 10251
rect 9689 10149 9723 10183
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 6837 10081 6871 10115
rect 9321 10081 9355 10115
rect 12173 10081 12207 10115
rect 3341 10013 3375 10047
rect 7205 10013 7239 10047
rect 7389 10013 7423 10047
rect 9873 10013 9907 10047
rect 10425 10013 10459 10047
rect 11437 10013 11471 10047
rect 11530 10013 11564 10047
rect 11902 10013 11936 10047
rect 12633 10013 12667 10047
rect 11713 9945 11747 9979
rect 11805 9945 11839 9979
rect 3157 9877 3191 9911
rect 10333 9877 10367 9911
rect 2881 9605 2915 9639
rect 4629 9605 4663 9639
rect 6009 9605 6043 9639
rect 9965 9605 9999 9639
rect 4721 9537 4755 9571
rect 5917 9537 5951 9571
rect 7481 9537 7515 9571
rect 7757 9537 7791 9571
rect 9689 9537 9723 9571
rect 9781 9537 9815 9571
rect 10793 9537 10827 9571
rect 11253 9537 11287 9571
rect 11805 9537 11839 9571
rect 12081 9537 12115 9571
rect 2605 9469 2639 9503
rect 8033 9469 8067 9503
rect 9505 9469 9539 9503
rect 9965 9469 9999 9503
rect 10977 9469 11011 9503
rect 11897 9469 11931 9503
rect 10885 9401 10919 9435
rect 4353 9333 4387 9367
rect 7389 9333 7423 9367
rect 10517 9333 10551 9367
rect 11069 9333 11103 9367
rect 11621 9333 11655 9367
rect 12081 9333 12115 9367
rect 8309 9129 8343 9163
rect 12265 9129 12299 9163
rect 4997 9061 5031 9095
rect 3249 8993 3283 9027
rect 4236 8993 4270 9027
rect 3525 8925 3559 8959
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 5457 8925 5491 8959
rect 7849 8925 7883 8959
rect 8217 8925 8251 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 12357 8925 12391 8959
rect 2973 8857 3007 8891
rect 5273 8857 5307 8891
rect 5733 8857 5767 8891
rect 1501 8789 1535 8823
rect 3433 8789 3467 8823
rect 4077 8789 4111 8823
rect 4353 8789 4387 8823
rect 4813 8789 4847 8823
rect 7205 8789 7239 8823
rect 7297 8789 7331 8823
rect 11437 8789 11471 8823
rect 3249 8585 3283 8619
rect 3341 8585 3375 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 2421 8517 2455 8551
rect 3525 8517 3559 8551
rect 3985 8517 4019 8551
rect 6377 8517 6411 8551
rect 12357 8517 12391 8551
rect 2329 8449 2363 8483
rect 2513 8449 2547 8483
rect 2605 8449 2639 8483
rect 2789 8449 2823 8483
rect 2881 8449 2915 8483
rect 2973 8449 3007 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 5917 8449 5951 8483
rect 6193 8449 6227 8483
rect 12081 8449 12115 8483
rect 12909 8381 12943 8415
rect 3893 8313 3927 8347
rect 12173 8313 12207 8347
rect 3525 8245 3559 8279
rect 7665 8245 7699 8279
rect 2605 8041 2639 8075
rect 3065 8041 3099 8075
rect 5549 8041 5583 8075
rect 12909 8041 12943 8075
rect 2237 7905 2271 7939
rect 9321 7905 9355 7939
rect 11437 7905 11471 7939
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 2789 7837 2823 7871
rect 2973 7837 3007 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 7021 7837 7055 7871
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 9689 7837 9723 7871
rect 11161 7837 11195 7871
rect 8953 7769 8987 7803
rect 9137 7769 9171 7803
rect 2237 7701 2271 7735
rect 8033 7701 8067 7735
rect 8401 7701 8435 7735
rect 9505 7701 9539 7735
rect 2697 7497 2731 7531
rect 5917 7497 5951 7531
rect 5733 7429 5767 7463
rect 8769 7429 8803 7463
rect 9505 7429 9539 7463
rect 2605 7361 2639 7395
rect 2789 7361 2823 7395
rect 6193 7361 6227 7395
rect 6561 7361 6595 7395
rect 9045 7361 9079 7395
rect 9229 7361 9263 7395
rect 11253 7361 11287 7395
rect 12173 7361 12207 7395
rect 11161 7293 11195 7327
rect 5365 7225 5399 7259
rect 5733 7157 5767 7191
rect 6009 7157 6043 7191
rect 6653 7157 6687 7191
rect 7297 7157 7331 7191
rect 10977 7157 11011 7191
rect 12265 7157 12299 7191
rect 1672 6953 1706 6987
rect 5812 6953 5846 6987
rect 8401 6953 8435 6987
rect 8585 6953 8619 6987
rect 9321 6953 9355 6987
rect 9965 6953 9999 6987
rect 10609 6953 10643 6987
rect 9137 6885 9171 6919
rect 5549 6817 5583 6851
rect 12909 6817 12943 6851
rect 1409 6749 1443 6783
rect 3433 6749 3467 6783
rect 4905 6749 4939 6783
rect 7573 6749 7607 6783
rect 7757 6749 7791 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 9689 6749 9723 6783
rect 10241 6749 10275 6783
rect 10885 6749 10919 6783
rect 11161 6749 11195 6783
rect 3341 6681 3375 6715
rect 4169 6681 4203 6715
rect 4353 6681 4387 6715
rect 5089 6681 5123 6715
rect 5273 6681 5307 6715
rect 5457 6681 5491 6715
rect 9321 6681 9355 6715
rect 10149 6681 10183 6715
rect 11437 6681 11471 6715
rect 3157 6613 3191 6647
rect 4537 6613 4571 6647
rect 4721 6613 4755 6647
rect 7297 6613 7331 6647
rect 8401 6613 8435 6647
rect 9781 6613 9815 6647
rect 9949 6613 9983 6647
rect 10609 6613 10643 6647
rect 10793 6613 10827 6647
rect 11069 6613 11103 6647
rect 3893 6409 3927 6443
rect 8585 6409 8619 6443
rect 9689 6409 9723 6443
rect 10333 6409 10367 6443
rect 4261 6341 4295 6375
rect 4629 6341 4663 6375
rect 9505 6341 9539 6375
rect 9873 6341 9907 6375
rect 9965 6341 9999 6375
rect 10149 6341 10183 6375
rect 4031 6307 4065 6341
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3525 6273 3559 6307
rect 4353 6273 4387 6307
rect 8217 6273 8251 6307
rect 8401 6273 8435 6307
rect 9597 6273 9631 6307
rect 12725 6273 12759 6307
rect 3341 6205 3375 6239
rect 3709 6205 3743 6239
rect 6101 6205 6135 6239
rect 9321 6205 9355 6239
rect 13001 6205 13035 6239
rect 2421 6069 2455 6103
rect 2789 6069 2823 6103
rect 4077 6069 4111 6103
rect 4353 5865 4387 5899
rect 5089 5865 5123 5899
rect 6469 5865 6503 5899
rect 3985 5797 4019 5831
rect 1501 5729 1535 5763
rect 1777 5729 1811 5763
rect 7941 5729 7975 5763
rect 8217 5729 8251 5763
rect 8309 5661 8343 5695
rect 4353 5593 4387 5627
rect 6377 5593 6411 5627
rect 8401 5593 8435 5627
rect 3249 5525 3283 5559
rect 4537 5525 4571 5559
rect 2789 5321 2823 5355
rect 4997 5321 5031 5355
rect 5365 5321 5399 5355
rect 5733 5321 5767 5355
rect 8769 5321 8803 5355
rect 10425 5321 10459 5355
rect 11345 5321 11379 5355
rect 2421 5253 2455 5287
rect 2973 5253 3007 5287
rect 3801 5253 3835 5287
rect 4169 5253 4203 5287
rect 5181 5253 5215 5287
rect 5549 5253 5583 5287
rect 8283 5253 8317 5287
rect 10517 5253 10551 5287
rect 10701 5253 10735 5287
rect 10977 5253 11011 5287
rect 11177 5253 11211 5287
rect 2145 5185 2179 5219
rect 3341 5185 3375 5219
rect 3985 5185 4019 5219
rect 5273 5185 5307 5219
rect 5825 5185 5859 5219
rect 7389 5185 7423 5219
rect 8401 5185 8435 5219
rect 8493 5185 8527 5219
rect 8585 5185 8619 5219
rect 9321 5185 9355 5219
rect 9781 5185 9815 5219
rect 10241 5185 10275 5219
rect 10425 5185 10459 5219
rect 11713 5185 11747 5219
rect 12173 5185 12207 5219
rect 8033 5117 8067 5151
rect 8125 5117 8159 5151
rect 2973 4981 3007 5015
rect 9229 4981 9263 5015
rect 9689 4981 9723 5015
rect 10885 4981 10919 5015
rect 11161 4981 11195 5015
rect 11529 4981 11563 5015
rect 12265 4981 12299 5015
rect 10701 4777 10735 4811
rect 2973 4641 3007 4675
rect 11437 4641 11471 4675
rect 1409 4573 1443 4607
rect 2697 4573 2731 4607
rect 10701 4573 10735 4607
rect 10885 4573 10919 4607
rect 11161 4573 11195 4607
rect 1593 4437 1627 4471
rect 12909 4437 12943 4471
rect 3341 4233 3375 4267
rect 4169 4233 4203 4267
rect 10241 4233 10275 4267
rect 10977 4233 11011 4267
rect 5641 4165 5675 4199
rect 7665 4165 7699 4199
rect 11161 4165 11195 4199
rect 2881 4097 2915 4131
rect 4537 4097 4571 4131
rect 4813 4097 4847 4131
rect 4905 4097 4939 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 8033 4097 8067 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 8677 4097 8711 4131
rect 8861 4097 8895 4131
rect 9413 4097 9447 4131
rect 10391 4097 10425 4131
rect 10885 4097 10919 4131
rect 11713 4097 11747 4131
rect 12357 4097 12391 4131
rect 12909 4097 12943 4131
rect 2237 4029 2271 4063
rect 3709 4029 3743 4063
rect 5825 4029 5859 4063
rect 6009 4029 6043 4063
rect 6745 4029 6779 4063
rect 10701 4029 10735 4063
rect 10793 4029 10827 4063
rect 11621 4029 11655 4063
rect 2605 3961 2639 3995
rect 4077 3961 4111 3995
rect 5273 3961 5307 3995
rect 7021 3961 7055 3995
rect 7113 3961 7147 3995
rect 7941 3961 7975 3995
rect 9137 3961 9171 3995
rect 11161 3961 11195 3995
rect 2697 3893 2731 3927
rect 3157 3893 3191 3927
rect 4629 3893 4663 3927
rect 5181 3893 5215 3927
rect 5917 3893 5951 3927
rect 8585 3893 8619 3927
rect 8861 3893 8895 3927
rect 9321 3893 9355 3927
rect 12081 3893 12115 3927
rect 1685 3689 1719 3723
rect 2329 3689 2363 3723
rect 2697 3689 2731 3723
rect 4537 3689 4571 3723
rect 5549 3689 5583 3723
rect 7021 3689 7055 3723
rect 7389 3689 7423 3723
rect 8953 3689 8987 3723
rect 10241 3689 10275 3723
rect 10977 3689 11011 3723
rect 12909 3689 12943 3723
rect 1961 3621 1995 3655
rect 2513 3621 2547 3655
rect 3525 3621 3559 3655
rect 5917 3621 5951 3655
rect 9413 3621 9447 3655
rect 4077 3553 4111 3587
rect 4169 3553 4203 3587
rect 5181 3553 5215 3587
rect 5733 3553 5767 3587
rect 6377 3553 6411 3587
rect 7113 3553 7147 3587
rect 8033 3553 8067 3587
rect 10517 3553 10551 3587
rect 11161 3553 11195 3587
rect 1409 3485 1443 3519
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4353 3485 4387 3519
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 5825 3485 5859 3519
rect 6101 3485 6135 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 7205 3485 7239 3519
rect 7606 3485 7640 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 8769 3485 8803 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 9487 3485 9521 3519
rect 9597 3485 9631 3519
rect 9690 3485 9724 3519
rect 9965 3485 9999 3519
rect 10062 3485 10096 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 10885 3485 10919 3519
rect 2973 3417 3007 3451
rect 6929 3417 6963 3451
rect 8493 3417 8527 3451
rect 9873 3417 9907 3451
rect 11437 3417 11471 3451
rect 1869 3349 1903 3383
rect 2329 3349 2363 3383
rect 2881 3349 2915 3383
rect 3341 3349 3375 3383
rect 7481 3349 7515 3383
rect 7665 3349 7699 3383
rect 8217 3349 8251 3383
rect 2973 3145 3007 3179
rect 3065 3145 3099 3179
rect 4445 3145 4479 3179
rect 5641 3145 5675 3179
rect 6929 3145 6963 3179
rect 7297 3145 7331 3179
rect 7941 3145 7975 3179
rect 8769 3145 8803 3179
rect 9689 3145 9723 3179
rect 12265 3145 12299 3179
rect 12541 3145 12575 3179
rect 3985 3077 4019 3111
rect 5273 3077 5307 3111
rect 6101 3077 6135 3111
rect 7573 3077 7607 3111
rect 8401 3077 8435 3111
rect 2513 3009 2547 3043
rect 3525 3009 3559 3043
rect 3877 3015 3911 3049
rect 4077 3009 4111 3043
rect 4261 3009 4295 3043
rect 4353 3009 4387 3043
rect 4905 3009 4939 3043
rect 5089 3009 5123 3043
rect 5365 3009 5399 3043
rect 5457 3009 5491 3043
rect 5917 3009 5951 3043
rect 6469 3009 6503 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 7757 3009 7791 3043
rect 8217 3009 8251 3043
rect 8493 3009 8527 3043
rect 8585 3009 8619 3043
rect 9137 3009 9171 3043
rect 9413 3009 9447 3043
rect 9505 3009 9539 3043
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 12449 3009 12483 3043
rect 13001 3009 13035 3043
rect 5733 2941 5767 2975
rect 6653 2941 6687 2975
rect 4537 2873 4571 2907
rect 9229 2873 9263 2907
rect 12817 2873 12851 2907
rect 2789 2805 2823 2839
rect 3433 2805 3467 2839
rect 3709 2805 3743 2839
rect 6469 2805 6503 2839
rect 1593 2601 1627 2635
rect 2789 2601 2823 2635
rect 4353 2601 4387 2635
rect 5917 2601 5951 2635
rect 8953 2601 8987 2635
rect 10425 2601 10459 2635
rect 12817 2601 12851 2635
rect 7297 2533 7331 2567
rect 11805 2465 11839 2499
rect 1409 2397 1443 2431
rect 2605 2397 2639 2431
rect 4169 2397 4203 2431
rect 5733 2397 5767 2431
rect 6745 2397 6779 2431
rect 6837 2397 6871 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 10609 2397 10643 2431
rect 11529 2397 11563 2431
rect 12909 2329 12943 2363
<< metal1 >>
rect 1104 14170 13340 14192
rect 1104 14118 3139 14170
rect 3191 14118 3203 14170
rect 3255 14118 3267 14170
rect 3319 14118 3331 14170
rect 3383 14118 3395 14170
rect 3447 14118 6198 14170
rect 6250 14118 6262 14170
rect 6314 14118 6326 14170
rect 6378 14118 6390 14170
rect 6442 14118 6454 14170
rect 6506 14118 9257 14170
rect 9309 14118 9321 14170
rect 9373 14118 9385 14170
rect 9437 14118 9449 14170
rect 9501 14118 9513 14170
rect 9565 14118 12316 14170
rect 12368 14118 12380 14170
rect 12432 14118 12444 14170
rect 12496 14118 12508 14170
rect 12560 14118 12572 14170
rect 12624 14118 13340 14170
rect 1104 14096 13340 14118
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 3660 14028 3893 14056
rect 3660 14016 3666 14028
rect 3881 14025 3893 14028
rect 3927 14025 3939 14059
rect 3881 14019 3939 14025
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10836 14028 11069 14056
rect 10836 14016 10842 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 12897 13991 12955 13997
rect 12897 13957 12909 13991
rect 12943 13988 12955 13991
rect 13262 13988 13268 14000
rect 12943 13960 13268 13988
rect 12943 13957 12955 13960
rect 12897 13951 12955 13957
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 12066 13744 12072 13796
rect 12124 13784 12130 13796
rect 12713 13787 12771 13793
rect 12713 13784 12725 13787
rect 12124 13756 12725 13784
rect 12124 13744 12130 13756
rect 12713 13753 12725 13756
rect 12759 13753 12771 13787
rect 12713 13747 12771 13753
rect 1104 13626 13340 13648
rect 1104 13574 2479 13626
rect 2531 13574 2543 13626
rect 2595 13574 2607 13626
rect 2659 13574 2671 13626
rect 2723 13574 2735 13626
rect 2787 13574 5538 13626
rect 5590 13574 5602 13626
rect 5654 13574 5666 13626
rect 5718 13574 5730 13626
rect 5782 13574 5794 13626
rect 5846 13574 8597 13626
rect 8649 13574 8661 13626
rect 8713 13574 8725 13626
rect 8777 13574 8789 13626
rect 8841 13574 8853 13626
rect 8905 13574 11656 13626
rect 11708 13574 11720 13626
rect 11772 13574 11784 13626
rect 11836 13574 11848 13626
rect 11900 13574 11912 13626
rect 11964 13574 13340 13626
rect 1104 13552 13340 13574
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6604 13348 6914 13376
rect 6604 13336 6610 13348
rect 6886 13240 6914 13348
rect 8018 13336 8024 13388
rect 8076 13376 8082 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 8076 13348 10241 13376
rect 8076 13336 8082 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7432 13280 7481 13308
rect 7432 13268 7438 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 8110 13268 8116 13320
rect 8168 13268 8174 13320
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9355 13280 9689 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 8956 13240 8984 13271
rect 6886 13212 8984 13240
rect 7466 13132 7472 13184
rect 7524 13132 7530 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7892 13144 7941 13172
rect 7892 13132 7898 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 9140 13172 9168 13271
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13209 10563 13243
rect 10505 13203 10563 13209
rect 8444 13144 9168 13172
rect 9861 13175 9919 13181
rect 8444 13132 8450 13144
rect 9861 13141 9873 13175
rect 9907 13172 9919 13175
rect 10520 13172 10548 13203
rect 9907 13144 10548 13172
rect 9907 13141 9919 13144
rect 9861 13135 9919 13141
rect 11974 13132 11980 13184
rect 12032 13132 12038 13184
rect 1104 13082 13340 13104
rect 1104 13030 3139 13082
rect 3191 13030 3203 13082
rect 3255 13030 3267 13082
rect 3319 13030 3331 13082
rect 3383 13030 3395 13082
rect 3447 13030 6198 13082
rect 6250 13030 6262 13082
rect 6314 13030 6326 13082
rect 6378 13030 6390 13082
rect 6442 13030 6454 13082
rect 6506 13030 9257 13082
rect 9309 13030 9321 13082
rect 9373 13030 9385 13082
rect 9437 13030 9449 13082
rect 9501 13030 9513 13082
rect 9565 13030 12316 13082
rect 12368 13030 12380 13082
rect 12432 13030 12444 13082
rect 12496 13030 12508 13082
rect 12560 13030 12572 13082
rect 12624 13030 13340 13082
rect 1104 13008 13340 13030
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7432 12940 9260 12968
rect 7432 12928 7438 12940
rect 6533 12903 6591 12909
rect 6533 12869 6545 12903
rect 6579 12900 6591 12903
rect 6638 12900 6644 12912
rect 6579 12872 6644 12900
rect 6579 12869 6591 12872
rect 6533 12863 6591 12869
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 6733 12903 6791 12909
rect 6733 12869 6745 12903
rect 6779 12869 6791 12903
rect 6733 12863 6791 12869
rect 7009 12903 7067 12909
rect 7009 12869 7021 12903
rect 7055 12900 7067 12903
rect 7282 12900 7288 12912
rect 7055 12872 7288 12900
rect 7055 12869 7067 12872
rect 7009 12863 7067 12869
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6135 12804 6408 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 5534 12724 5540 12776
rect 5592 12764 5598 12776
rect 5644 12764 5672 12795
rect 5592 12736 5672 12764
rect 5721 12767 5779 12773
rect 5592 12724 5598 12736
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 5902 12764 5908 12776
rect 5767 12736 5908 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6380 12705 6408 12804
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 6748 12764 6776 12863
rect 7282 12860 7288 12872
rect 7340 12860 7346 12912
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 7392 12832 7420 12928
rect 8018 12900 8024 12912
rect 7484 12872 8024 12900
rect 7484 12841 7512 12872
rect 8018 12860 8024 12872
rect 8076 12860 8082 12912
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 7239 12804 7420 12832
rect 7469 12835 7527 12841
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 6604 12736 6776 12764
rect 7745 12767 7803 12773
rect 6604 12724 6610 12736
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 7834 12764 7840 12776
rect 7791 12736 7840 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 9232 12773 9260 12940
rect 11606 12928 11612 12980
rect 11664 12928 11670 12980
rect 10704 12872 12112 12900
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 10704 12841 10732 12872
rect 12084 12844 12112 12872
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9732 12804 9781 12832
rect 9732 12792 9738 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 11422 12792 11428 12844
rect 11480 12832 11486 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11480 12804 11713 12832
rect 11480 12792 11486 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 12066 12792 12072 12844
rect 12124 12792 12130 12844
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9263 12736 9505 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 9493 12733 9505 12736
rect 9539 12764 9551 12767
rect 10134 12764 10140 12776
rect 9539 12736 10140 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 6365 12699 6423 12705
rect 6365 12665 6377 12699
rect 6411 12665 6423 12699
rect 6365 12659 6423 12665
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 9858 12696 9864 12708
rect 9631 12668 9864 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 9858 12656 9864 12668
rect 9916 12696 9922 12708
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 9916 12668 10609 12696
rect 9916 12656 9922 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 5905 12631 5963 12637
rect 5905 12597 5917 12631
rect 5951 12628 5963 12631
rect 5994 12628 6000 12640
rect 5951 12600 6000 12628
rect 5951 12597 5963 12600
rect 5905 12591 5963 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 7190 12628 7196 12640
rect 6595 12600 7196 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7374 12588 7380 12640
rect 7432 12588 7438 12640
rect 9953 12631 10011 12637
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10318 12628 10324 12640
rect 9999 12600 10324 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 1104 12538 13340 12560
rect 1104 12486 2479 12538
rect 2531 12486 2543 12538
rect 2595 12486 2607 12538
rect 2659 12486 2671 12538
rect 2723 12486 2735 12538
rect 2787 12486 5538 12538
rect 5590 12486 5602 12538
rect 5654 12486 5666 12538
rect 5718 12486 5730 12538
rect 5782 12486 5794 12538
rect 5846 12486 8597 12538
rect 8649 12486 8661 12538
rect 8713 12486 8725 12538
rect 8777 12486 8789 12538
rect 8841 12486 8853 12538
rect 8905 12486 11656 12538
rect 11708 12486 11720 12538
rect 11772 12486 11784 12538
rect 11836 12486 11848 12538
rect 11900 12486 11912 12538
rect 11964 12486 13340 12538
rect 1104 12464 13340 12486
rect 7377 12427 7435 12433
rect 7377 12393 7389 12427
rect 7423 12424 7435 12427
rect 7466 12424 7472 12436
rect 7423 12396 7472 12424
rect 7423 12393 7435 12396
rect 7377 12387 7435 12393
rect 7466 12384 7472 12396
rect 7524 12424 7530 12436
rect 7524 12396 8156 12424
rect 7524 12384 7530 12396
rect 7561 12359 7619 12365
rect 6472 12328 7512 12356
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 6472 12288 6500 12328
rect 5132 12260 6500 12288
rect 5132 12248 5138 12260
rect 6546 12248 6552 12300
rect 6604 12248 6610 12300
rect 6564 12220 6592 12248
rect 6730 12220 6736 12232
rect 6564 12192 6736 12220
rect 6730 12180 6736 12192
rect 6788 12220 6794 12232
rect 7484 12220 7512 12328
rect 7561 12325 7573 12359
rect 7607 12325 7619 12359
rect 7561 12319 7619 12325
rect 7576 12288 7604 12319
rect 8128 12297 8156 12396
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8536 12396 8585 12424
rect 8536 12384 8542 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 9674 12384 9680 12436
rect 9732 12384 9738 12436
rect 10410 12424 10416 12436
rect 9784 12396 10416 12424
rect 8386 12316 8392 12368
rect 8444 12316 8450 12368
rect 9784 12365 9812 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 11974 12424 11980 12436
rect 11931 12396 11980 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 9769 12359 9827 12365
rect 9769 12325 9781 12359
rect 9815 12325 9827 12359
rect 11900 12356 11928 12387
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 9769 12319 9827 12325
rect 9876 12328 11928 12356
rect 8113 12291 8171 12297
rect 7576 12260 7880 12288
rect 7742 12220 7748 12232
rect 6788 12192 7236 12220
rect 7484 12192 7748 12220
rect 6788 12180 6794 12192
rect 5353 12155 5411 12161
rect 5353 12121 5365 12155
rect 5399 12121 5411 12155
rect 5353 12115 5411 12121
rect 5368 12084 5396 12115
rect 5902 12112 5908 12164
rect 5960 12112 5966 12164
rect 7208 12161 7236 12192
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 7193 12155 7251 12161
rect 7193 12121 7205 12155
rect 7239 12121 7251 12155
rect 7193 12115 7251 12121
rect 7374 12112 7380 12164
rect 7432 12161 7438 12164
rect 7432 12155 7451 12161
rect 7439 12121 7451 12155
rect 7852 12152 7880 12260
rect 8113 12257 8125 12291
rect 8159 12257 8171 12291
rect 9876 12288 9904 12328
rect 8113 12251 8171 12257
rect 8404 12260 9904 12288
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12220 8079 12223
rect 8404 12220 8432 12260
rect 10331 12233 10389 12239
rect 8067 12192 8432 12220
rect 8481 12223 8539 12229
rect 8067 12189 8079 12192
rect 8021 12183 8079 12189
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8110 12152 8116 12164
rect 7852 12124 8116 12152
rect 7432 12115 7451 12121
rect 7432 12112 7438 12115
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 8386 12112 8392 12164
rect 8444 12152 8450 12164
rect 8496 12152 8524 12183
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 8444 12124 8524 12152
rect 8444 12112 8450 12124
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 9088 12124 9321 12152
rect 9088 12112 9094 12124
rect 9309 12121 9321 12124
rect 9355 12121 9367 12155
rect 9309 12115 9367 12121
rect 9401 12155 9459 12161
rect 9401 12121 9413 12155
rect 9447 12121 9459 12155
rect 9508 12152 9536 12183
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10134 12229 10140 12232
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9916 12192 9965 12220
rect 9916 12180 9922 12192
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10118 12223 10140 12229
rect 10118 12189 10130 12223
rect 10118 12183 10140 12189
rect 10134 12180 10140 12183
rect 10192 12180 10198 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10331 12199 10343 12233
rect 10377 12230 10389 12233
rect 10428 12230 10456 12328
rect 10377 12202 10456 12230
rect 11977 12223 12035 12229
rect 10377 12199 10389 12202
rect 10331 12193 10389 12199
rect 10229 12183 10287 12189
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12066 12220 12072 12232
rect 12023 12192 12072 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 9508 12124 9996 12152
rect 9401 12115 9459 12121
rect 5994 12084 6000 12096
rect 5368 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6825 12087 6883 12093
rect 6825 12053 6837 12087
rect 6871 12084 6883 12087
rect 7098 12084 7104 12096
rect 6871 12056 7104 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7098 12044 7104 12056
rect 7156 12084 7162 12096
rect 9416 12084 9444 12115
rect 9968 12096 9996 12124
rect 9628 12084 9634 12096
rect 7156 12056 9634 12084
rect 7156 12044 7162 12056
rect 9628 12044 9634 12056
rect 9686 12044 9692 12096
rect 9950 12044 9956 12096
rect 10008 12044 10014 12096
rect 10244 12084 10272 12183
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 10318 12084 10324 12096
rect 10244 12056 10324 12084
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 11514 12044 11520 12096
rect 11572 12044 11578 12096
rect 1104 11994 13340 12016
rect 1104 11942 3139 11994
rect 3191 11942 3203 11994
rect 3255 11942 3267 11994
rect 3319 11942 3331 11994
rect 3383 11942 3395 11994
rect 3447 11942 6198 11994
rect 6250 11942 6262 11994
rect 6314 11942 6326 11994
rect 6378 11942 6390 11994
rect 6442 11942 6454 11994
rect 6506 11942 9257 11994
rect 9309 11942 9321 11994
rect 9373 11942 9385 11994
rect 9437 11942 9449 11994
rect 9501 11942 9513 11994
rect 9565 11942 12316 11994
rect 12368 11942 12380 11994
rect 12432 11942 12444 11994
rect 12496 11942 12508 11994
rect 12560 11942 12572 11994
rect 12624 11942 13340 11994
rect 1104 11920 13340 11942
rect 7009 11883 7067 11889
rect 6656 11852 6960 11880
rect 6656 11821 6684 11852
rect 6641 11815 6699 11821
rect 6641 11781 6653 11815
rect 6687 11781 6699 11815
rect 6841 11815 6899 11821
rect 6841 11812 6853 11815
rect 6641 11775 6699 11781
rect 6748 11784 6853 11812
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 5902 11744 5908 11756
rect 4847 11716 5908 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 6748 11744 6776 11784
rect 6841 11781 6853 11784
rect 6887 11781 6899 11815
rect 6841 11775 6899 11781
rect 6604 11716 6776 11744
rect 6932 11744 6960 11852
rect 7009 11849 7021 11883
rect 7055 11849 7067 11883
rect 7009 11843 7067 11849
rect 7024 11812 7052 11843
rect 7190 11840 7196 11892
rect 7248 11840 7254 11892
rect 7282 11840 7288 11892
rect 7340 11840 7346 11892
rect 9490 11840 9496 11892
rect 9548 11840 9554 11892
rect 10042 11880 10048 11892
rect 9876 11852 10048 11880
rect 7300 11812 7328 11840
rect 7024 11784 7328 11812
rect 7098 11744 7104 11756
rect 6932 11716 7104 11744
rect 6604 11704 6610 11716
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 7300 11753 7328 11784
rect 9508 11753 9536 11840
rect 9769 11815 9827 11821
rect 9769 11781 9781 11815
rect 9815 11812 9827 11815
rect 9876 11812 9904 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 10284 11852 11100 11880
rect 10284 11840 10290 11852
rect 9815 11784 9904 11812
rect 10336 11784 11008 11812
rect 9815 11781 9827 11784
rect 9769 11775 9827 11781
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 8386 11676 8392 11688
rect 5592 11648 8392 11676
rect 5592 11636 5598 11648
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 9122 11636 9128 11688
rect 9180 11636 9186 11688
rect 9416 11676 9444 11707
rect 9582 11704 9588 11756
rect 9640 11704 9646 11756
rect 9950 11704 9956 11756
rect 10008 11744 10014 11756
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 10008 11716 10057 11744
rect 10008 11704 10014 11716
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 10060 11676 10088 11707
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10336 11744 10364 11784
rect 10980 11756 11008 11784
rect 10192 11716 10364 11744
rect 10192 11704 10198 11716
rect 10410 11704 10416 11756
rect 10468 11704 10474 11756
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 11072 11753 11100 11852
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11103 11716 11713 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11992 11744 12020 11840
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11992 11716 12173 11744
rect 11701 11707 11759 11713
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 11333 11679 11391 11685
rect 9416 11648 9536 11676
rect 9140 11608 9168 11636
rect 9508 11608 9536 11648
rect 10060 11648 11192 11676
rect 10060 11608 10088 11648
rect 9140 11580 9444 11608
rect 9508 11580 10088 11608
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4396 11512 4629 11540
rect 4396 11500 4402 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7190 11540 7196 11552
rect 6871 11512 7196 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8352 11512 9229 11540
rect 8352 11500 8358 11512
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9416 11540 9444 11580
rect 11164 11552 11192 11648
rect 11333 11645 11345 11679
rect 11379 11676 11391 11679
rect 11514 11676 11520 11688
rect 11379 11648 11520 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11624 11608 11652 11639
rect 11440 11580 11652 11608
rect 11440 11552 11468 11580
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9416 11512 9873 11540
rect 9217 11503 9275 11509
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 9861 11503 9919 11509
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10686 11540 10692 11552
rect 10367 11512 10692 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11146 11500 11152 11552
rect 11204 11500 11210 11552
rect 11238 11500 11244 11552
rect 11296 11500 11302 11552
rect 11422 11500 11428 11552
rect 11480 11500 11486 11552
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12250 11500 12256 11552
rect 12308 11500 12314 11552
rect 1104 11450 13340 11472
rect 1104 11398 2479 11450
rect 2531 11398 2543 11450
rect 2595 11398 2607 11450
rect 2659 11398 2671 11450
rect 2723 11398 2735 11450
rect 2787 11398 5538 11450
rect 5590 11398 5602 11450
rect 5654 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 8597 11450
rect 8649 11398 8661 11450
rect 8713 11398 8725 11450
rect 8777 11398 8789 11450
rect 8841 11398 8853 11450
rect 8905 11398 11656 11450
rect 11708 11398 11720 11450
rect 11772 11398 11784 11450
rect 11836 11398 11848 11450
rect 11900 11398 11912 11450
rect 11964 11398 13340 11450
rect 1104 11376 13340 11398
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 5994 11336 6000 11348
rect 4120 11308 6000 11336
rect 4120 11296 4126 11308
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6696 11308 6837 11336
rect 6696 11296 6702 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 9030 11296 9036 11348
rect 9088 11296 9094 11348
rect 10686 11296 10692 11348
rect 10744 11296 10750 11348
rect 11146 11296 11152 11348
rect 11204 11296 11210 11348
rect 12250 11296 12256 11348
rect 12308 11296 12314 11348
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 8113 11271 8171 11277
rect 8113 11268 8125 11271
rect 6788 11240 8125 11268
rect 6788 11228 6794 11240
rect 8113 11237 8125 11240
rect 8159 11237 8171 11271
rect 10042 11268 10048 11280
rect 8113 11231 8171 11237
rect 9324 11240 10048 11268
rect 3789 11203 3847 11209
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 6181 11203 6239 11209
rect 3835 11172 5120 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 5092 11144 5120 11172
rect 6181 11169 6193 11203
rect 6227 11200 6239 11203
rect 6546 11200 6552 11212
rect 6227 11172 6552 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 9324 11200 9352 11240
rect 10042 11228 10048 11240
rect 10100 11268 10106 11280
rect 10704 11268 10732 11296
rect 11422 11268 11428 11280
rect 10100 11240 10732 11268
rect 11256 11240 11428 11268
rect 10100 11228 10106 11240
rect 10502 11200 10508 11212
rect 7147 11172 7420 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 7392 11144 7420 11172
rect 9232 11172 9352 11200
rect 9646 11172 10508 11200
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4338 11064 4344 11076
rect 4111 11036 4344 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 4706 11024 4712 11076
rect 4764 11024 4770 11076
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 6104 11064 6132 11095
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7282 11092 7288 11144
rect 7340 11092 7346 11144
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 9232 11141 9260 11172
rect 9646 11151 9674 11172
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 9595 11145 9674 11151
rect 9217 11135 9275 11141
rect 7484 11104 9168 11132
rect 7208 11064 7236 11092
rect 7484 11064 7512 11104
rect 5859 11036 7512 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 8294 11024 8300 11076
rect 8352 11024 8358 11076
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 8444 11036 8493 11064
rect 8444 11024 8450 11036
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 9140 11064 9168 11104
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 9595 11111 9607 11145
rect 9641 11114 9674 11145
rect 9641 11111 9653 11114
rect 9595 11105 9653 11111
rect 9493 11095 9551 11101
rect 9324 11064 9352 11095
rect 9140 11036 9352 11064
rect 9508 11064 9536 11095
rect 10410 11092 10416 11144
rect 10468 11092 10474 11144
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11256 11141 11284 11240
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 12268 11200 12296 11296
rect 11348 11172 11836 11200
rect 11348 11144 11376 11172
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 11204 11104 11253 11132
rect 11204 11092 11210 11104
rect 11241 11101 11253 11104
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 11514 11132 11520 11144
rect 11471 11104 11520 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 9582 11064 9588 11076
rect 9508 11036 9588 11064
rect 8481 11027 8539 11033
rect 6457 10999 6515 11005
rect 6457 10965 6469 10999
rect 6503 10996 6515 10999
rect 6638 10996 6644 11008
rect 6503 10968 6644 10996
rect 6503 10965 6515 10968
rect 6457 10959 6515 10965
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 9324 10996 9352 11036
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 9950 10996 9956 11008
rect 9324 10968 9956 10996
rect 9950 10956 9956 10968
rect 10008 10996 10014 11008
rect 10428 10996 10456 11092
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 11072 11036 11713 11064
rect 11072 11008 11100 11036
rect 11701 11033 11713 11036
rect 11747 11033 11759 11067
rect 11808 11064 11836 11172
rect 11992 11172 12296 11200
rect 11992 11141 12020 11172
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12084 11064 12112 11092
rect 11808 11036 12112 11064
rect 11701 11027 11759 11033
rect 10008 10968 10456 10996
rect 10008 10956 10014 10968
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 11514 10956 11520 11008
rect 11572 10956 11578 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12360 10996 12388 11095
rect 12124 10968 12388 10996
rect 12124 10956 12130 10968
rect 1104 10906 13340 10928
rect 1104 10854 3139 10906
rect 3191 10854 3203 10906
rect 3255 10854 3267 10906
rect 3319 10854 3331 10906
rect 3383 10854 3395 10906
rect 3447 10854 6198 10906
rect 6250 10854 6262 10906
rect 6314 10854 6326 10906
rect 6378 10854 6390 10906
rect 6442 10854 6454 10906
rect 6506 10854 9257 10906
rect 9309 10854 9321 10906
rect 9373 10854 9385 10906
rect 9437 10854 9449 10906
rect 9501 10854 9513 10906
rect 9565 10854 12316 10906
rect 12368 10854 12380 10906
rect 12432 10854 12444 10906
rect 12496 10854 12508 10906
rect 12560 10854 12572 10906
rect 12624 10854 13340 10906
rect 1104 10832 13340 10854
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 5960 10764 6377 10792
rect 5960 10752 5966 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 6365 10755 6423 10761
rect 6564 10764 8033 10792
rect 6564 10724 6592 10764
rect 8021 10761 8033 10764
rect 8067 10761 8079 10795
rect 10226 10792 10232 10804
rect 8021 10755 8079 10761
rect 9692 10764 10232 10792
rect 5920 10696 6592 10724
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 4798 10656 4804 10668
rect 4663 10628 4804 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 4798 10616 4804 10628
rect 4856 10656 4862 10668
rect 5442 10656 5448 10668
rect 4856 10628 5448 10656
rect 4856 10616 4862 10628
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5920 10665 5948 10696
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6696 10696 6837 10724
rect 6696 10684 6702 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 7024 10696 8156 10724
rect 7024 10668 7052 10696
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10625 6147 10659
rect 6089 10619 6147 10625
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10656 6239 10659
rect 6227 10628 6592 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 5902 10412 5908 10464
rect 5960 10412 5966 10464
rect 6104 10452 6132 10619
rect 6564 10600 6592 10628
rect 7006 10616 7012 10668
rect 7064 10616 7070 10668
rect 8128 10665 8156 10696
rect 8386 10684 8392 10736
rect 8444 10724 8450 10736
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 8444 10696 9597 10724
rect 8444 10684 8450 10696
rect 9585 10693 9597 10696
rect 9631 10693 9643 10727
rect 9585 10687 9643 10693
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7883 10628 7941 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 8294 10656 8300 10668
rect 8251 10628 8300 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 9692 10656 9720 10764
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10686 10752 10692 10804
rect 10744 10752 10750 10804
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11885 10795 11943 10801
rect 11020 10764 11652 10792
rect 11020 10752 11026 10764
rect 11624 10724 11652 10764
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11974 10792 11980 10804
rect 11931 10764 11980 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12618 10724 12624 10736
rect 9968 10696 11560 10724
rect 11624 10696 12624 10724
rect 8527 10628 9720 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 9766 10616 9772 10668
rect 9824 10616 9830 10668
rect 9968 10665 9996 10696
rect 11532 10668 11560 10696
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 7374 10588 7380 10600
rect 7331 10560 7380 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 10060 10588 10088 10619
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 10827 10628 11192 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 10873 10591 10931 10597
rect 8128 10560 10824 10588
rect 6457 10523 6515 10529
rect 6457 10489 6469 10523
rect 6503 10520 6515 10523
rect 6730 10520 6736 10532
rect 6503 10492 6736 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 8128 10452 8156 10560
rect 9861 10523 9919 10529
rect 9861 10489 9873 10523
rect 9907 10520 9919 10523
rect 10594 10520 10600 10532
rect 9907 10492 10600 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10796 10520 10824 10560
rect 10873 10557 10885 10591
rect 10919 10588 10931 10591
rect 10962 10588 10968 10600
rect 10919 10560 10968 10588
rect 10919 10557 10931 10560
rect 10873 10551 10931 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11054 10520 11060 10532
rect 10796 10492 11060 10520
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11164 10529 11192 10628
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12250 10656 12256 10668
rect 12124 10628 12256 10656
rect 12124 10616 12130 10628
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 12342 10616 12348 10668
rect 12400 10656 12406 10668
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12400 10628 12725 10656
rect 12400 10616 12406 10628
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12713 10619 12771 10625
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11606 10588 11612 10600
rect 11480 10560 11612 10588
rect 11480 10548 11486 10560
rect 11606 10548 11612 10560
rect 11664 10588 11670 10600
rect 11664 10560 12112 10588
rect 11664 10548 11670 10560
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10489 11207 10523
rect 11149 10483 11207 10489
rect 11333 10523 11391 10529
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 11514 10520 11520 10532
rect 11379 10492 11520 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 6104 10424 8156 10452
rect 8205 10455 8263 10461
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 8386 10452 8392 10464
rect 8251 10424 8392 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9640 10424 10333 10452
rect 9640 10412 9646 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 11164 10452 11192 10483
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 12084 10529 12112 10560
rect 12986 10548 12992 10600
rect 13044 10548 13050 10600
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 11020 10424 11192 10452
rect 11885 10455 11943 10461
rect 11020 10412 11026 10424
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 11974 10452 11980 10464
rect 11931 10424 11980 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 1104 10362 13340 10384
rect 1104 10310 2479 10362
rect 2531 10310 2543 10362
rect 2595 10310 2607 10362
rect 2659 10310 2671 10362
rect 2723 10310 2735 10362
rect 2787 10310 5538 10362
rect 5590 10310 5602 10362
rect 5654 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 8597 10362
rect 8649 10310 8661 10362
rect 8713 10310 8725 10362
rect 8777 10310 8789 10362
rect 8841 10310 8853 10362
rect 8905 10310 11656 10362
rect 11708 10310 11720 10362
rect 11772 10310 11784 10362
rect 11836 10310 11848 10362
rect 11900 10310 11912 10362
rect 11964 10310 13340 10362
rect 1104 10288 13340 10310
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6604 10220 7021 10248
rect 6604 10208 6610 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 9766 10208 9772 10260
rect 9824 10208 9830 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 10502 10208 10508 10260
rect 10560 10208 10566 10260
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10652 10220 10885 10248
rect 10652 10208 10658 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11698 10248 11704 10260
rect 11020 10220 11704 10248
rect 11020 10208 11026 10220
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 12158 10248 12164 10260
rect 12115 10220 12164 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10217 12403 10251
rect 12345 10211 12403 10217
rect 9677 10183 9735 10189
rect 9677 10149 9689 10183
rect 9723 10180 9735 10183
rect 9968 10180 9996 10208
rect 9723 10152 9996 10180
rect 9723 10149 9735 10152
rect 9677 10143 9735 10149
rect 10410 10140 10416 10192
rect 10468 10140 10474 10192
rect 5074 10072 5080 10124
rect 5132 10072 5138 10124
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5902 10112 5908 10124
rect 5399 10084 5908 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 9309 10115 9367 10121
rect 6871 10084 7420 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7392 10056 7420 10084
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 10428 10112 10456 10140
rect 11054 10112 11060 10124
rect 9355 10084 11060 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 3602 10044 3608 10056
rect 3375 10016 3608 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 7116 10016 7205 10044
rect 5902 9936 5908 9988
rect 5960 9936 5966 9988
rect 7116 9920 7144 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7374 10004 7380 10056
rect 7432 10004 7438 10056
rect 9876 10053 9904 10084
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11606 10072 11612 10124
rect 11664 10072 11670 10124
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 12032 10084 12173 10112
rect 12032 10072 12038 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9861 10007 9919 10013
rect 10336 10016 10425 10044
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3145 9911 3203 9917
rect 3145 9908 3157 9911
rect 3016 9880 3157 9908
rect 3016 9868 3022 9880
rect 3145 9877 3157 9880
rect 3191 9877 3203 9911
rect 3145 9871 3203 9877
rect 7098 9868 7104 9920
rect 7156 9868 7162 9920
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10336 9917 10364 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11296 10016 11437 10044
rect 11296 10004 11302 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11624 10044 11652 10072
rect 11890 10047 11948 10053
rect 11890 10046 11902 10047
rect 11808 10044 11902 10046
rect 11624 10018 11902 10044
rect 11624 10016 11836 10018
rect 11890 10013 11902 10018
rect 11936 10013 11948 10047
rect 11890 10007 11948 10013
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9945 11759 9979
rect 11701 9939 11759 9945
rect 11793 9979 11851 9985
rect 11793 9945 11805 9979
rect 11839 9945 11851 9979
rect 12360 9976 12388 10211
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 11793 9939 11851 9945
rect 11992 9948 12388 9976
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10008 9880 10333 9908
rect 10008 9868 10014 9880
rect 10321 9877 10333 9880
rect 10367 9877 10379 9911
rect 10321 9871 10379 9877
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 11716 9908 11744 9939
rect 11480 9880 11744 9908
rect 11808 9908 11836 9939
rect 11992 9920 12020 9948
rect 11882 9908 11888 9920
rect 11808 9880 11888 9908
rect 11480 9868 11486 9880
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 11974 9868 11980 9920
rect 12032 9868 12038 9920
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 12342 9908 12348 9920
rect 12124 9880 12348 9908
rect 12124 9868 12130 9880
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 1104 9818 13340 9840
rect 1104 9766 3139 9818
rect 3191 9766 3203 9818
rect 3255 9766 3267 9818
rect 3319 9766 3331 9818
rect 3383 9766 3395 9818
rect 3447 9766 6198 9818
rect 6250 9766 6262 9818
rect 6314 9766 6326 9818
rect 6378 9766 6390 9818
rect 6442 9766 6454 9818
rect 6506 9766 9257 9818
rect 9309 9766 9321 9818
rect 9373 9766 9385 9818
rect 9437 9766 9449 9818
rect 9501 9766 9513 9818
rect 9565 9766 12316 9818
rect 12368 9766 12380 9818
rect 12432 9766 12444 9818
rect 12496 9766 12508 9818
rect 12560 9766 12572 9818
rect 12624 9766 13340 9818
rect 1104 9744 13340 9766
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 4856 9676 5856 9704
rect 4856 9664 4862 9676
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 2958 9636 2964 9648
rect 2915 9608 2964 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 4094 9608 4629 9636
rect 4617 9605 4629 9608
rect 4663 9605 4675 9639
rect 4617 9599 4675 9605
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4264 9540 4721 9568
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9469 2651 9503
rect 2593 9463 2651 9469
rect 2608 9364 2636 9463
rect 3234 9364 3240 9376
rect 2608 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 4264 9364 4292 9540
rect 4709 9537 4721 9540
rect 4755 9537 4767 9571
rect 5828 9568 5856 9676
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 5960 9676 6040 9704
rect 5960 9664 5966 9676
rect 6012 9645 6040 9676
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 10502 9704 10508 9716
rect 7432 9676 10508 9704
rect 7432 9664 7438 9676
rect 5997 9639 6055 9645
rect 5997 9605 6009 9639
rect 6043 9605 6055 9639
rect 5997 9599 6055 9605
rect 8478 9596 8484 9648
rect 8536 9596 8542 9648
rect 5905 9571 5963 9577
rect 5905 9568 5917 9571
rect 5828 9540 5917 9568
rect 4709 9531 4767 9537
rect 5905 9537 5917 9540
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 4724 9500 4752 9531
rect 7484 9500 7512 9531
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 9692 9577 9720 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11514 9664 11520 9716
rect 11572 9664 11578 9716
rect 9953 9639 10011 9645
rect 9953 9605 9965 9639
rect 9999 9636 10011 9639
rect 11532 9636 11560 9664
rect 9999 9608 11560 9636
rect 9999 9605 10011 9608
rect 9953 9599 10011 9605
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9537 9735 9571
rect 9677 9531 9735 9537
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 9876 9540 10793 9568
rect 4724 9472 7512 9500
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8386 9500 8392 9512
rect 8067 9472 8392 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9500 9551 9503
rect 9876 9500 9904 9540
rect 10781 9537 10793 9540
rect 10827 9568 10839 9571
rect 10870 9568 10876 9580
rect 10827 9540 10876 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11698 9568 11704 9580
rect 11287 9540 11704 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11698 9528 11704 9540
rect 11756 9568 11762 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11756 9540 11805 9568
rect 11756 9528 11762 9540
rect 11793 9537 11805 9540
rect 11839 9568 11851 9571
rect 11974 9568 11980 9580
rect 11839 9540 11980 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12066 9528 12072 9580
rect 12124 9528 12130 9580
rect 9539 9472 9904 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9950 9460 9956 9512
rect 10008 9460 10014 9512
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11330 9500 11336 9512
rect 11011 9472 11336 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11330 9460 11336 9472
rect 11388 9500 11394 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11388 9472 11897 9500
rect 11388 9460 11394 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 10873 9435 10931 9441
rect 10873 9401 10885 9435
rect 10919 9432 10931 9435
rect 11146 9432 11152 9444
rect 10919 9404 11152 9432
rect 10919 9401 10931 9404
rect 10873 9395 10931 9401
rect 11146 9392 11152 9404
rect 11204 9432 11210 9444
rect 12084 9432 12112 9528
rect 11204 9404 12112 9432
rect 11204 9392 11210 9404
rect 3568 9336 4292 9364
rect 3568 9324 3574 9336
rect 4338 9324 4344 9376
rect 4396 9324 4402 9376
rect 7374 9324 7380 9376
rect 7432 9324 7438 9376
rect 10502 9324 10508 9376
rect 10560 9324 10566 9376
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11422 9364 11428 9376
rect 11112 9336 11428 9364
rect 11112 9324 11118 9336
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11572 9336 11621 9364
rect 11572 9324 11578 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11756 9336 12081 9364
rect 11756 9324 11762 9336
rect 12069 9333 12081 9336
rect 12115 9364 12127 9367
rect 13078 9364 13084 9376
rect 12115 9336 13084 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 1104 9274 13340 9296
rect 1104 9222 2479 9274
rect 2531 9222 2543 9274
rect 2595 9222 2607 9274
rect 2659 9222 2671 9274
rect 2723 9222 2735 9274
rect 2787 9222 5538 9274
rect 5590 9222 5602 9274
rect 5654 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 8597 9274
rect 8649 9222 8661 9274
rect 8713 9222 8725 9274
rect 8777 9222 8789 9274
rect 8841 9222 8853 9274
rect 8905 9222 11656 9274
rect 11708 9222 11720 9274
rect 11772 9222 11784 9274
rect 11836 9222 11848 9274
rect 11900 9222 11912 9274
rect 11964 9222 13340 9274
rect 1104 9200 13340 9222
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 5074 9160 5080 9172
rect 3292 9132 5080 9160
rect 3292 9120 3298 9132
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 7374 9120 7380 9172
rect 7432 9120 7438 9172
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8478 9160 8484 9172
rect 8343 9132 8484 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 12253 9163 12311 9169
rect 12253 9160 12265 9163
rect 12216 9132 12265 9160
rect 12216 9120 12222 9132
rect 12253 9129 12265 9132
rect 12299 9129 12311 9163
rect 12253 9123 12311 9129
rect 3252 9033 3280 9120
rect 4985 9095 5043 9101
rect 4985 9092 4997 9095
rect 4448 9064 4997 9092
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 8993 3295 9027
rect 3237 8987 3295 8993
rect 4224 9027 4282 9033
rect 4224 8993 4236 9027
rect 4270 9024 4282 9027
rect 4338 9024 4344 9036
rect 4270 8996 4344 9024
rect 4270 8993 4282 8996
rect 4224 8987 4282 8993
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 4448 8965 4476 9064
rect 4985 9061 4997 9064
rect 5031 9092 5043 9095
rect 7392 9092 7420 9120
rect 11514 9092 11520 9104
rect 5031 9064 5396 9092
rect 5031 9061 5043 9064
rect 4985 9055 5043 9061
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 4755 8928 5304 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 2530 8860 2636 8888
rect 1486 8780 1492 8832
rect 1544 8780 1550 8832
rect 2608 8820 2636 8860
rect 2958 8848 2964 8900
rect 3016 8848 3022 8900
rect 3528 8832 3556 8919
rect 5276 8897 5304 8928
rect 5261 8891 5319 8897
rect 5261 8857 5273 8891
rect 5307 8857 5319 8891
rect 5368 8888 5396 9064
rect 6840 9064 7420 9092
rect 11348 9064 11520 9092
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 6840 8942 6868 9064
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 11348 9024 11376 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 12176 9024 12204 9120
rect 7156 8996 11376 9024
rect 7156 8984 7162 8996
rect 11348 8965 11376 8996
rect 11532 8996 12204 9024
rect 11532 8965 11560 8996
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8925 7895 8959
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 7837 8919 7895 8925
rect 8128 8928 8217 8956
rect 5626 8888 5632 8900
rect 5368 8860 5632 8888
rect 5261 8851 5319 8857
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 2608 8792 3433 8820
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3510 8780 3516 8832
rect 3568 8780 3574 8832
rect 4062 8780 4068 8832
rect 4120 8780 4126 8832
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4488 8792 4813 8820
rect 4488 8780 4494 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 5276 8820 5304 8851
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 5718 8848 5724 8900
rect 5776 8848 5782 8900
rect 7852 8888 7880 8919
rect 7208 8860 7880 8888
rect 7208 8829 7236 8860
rect 8128 8832 8156 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 12216 8928 12357 8956
rect 12216 8916 12222 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 5276 8792 7205 8820
rect 4801 8783 4859 8789
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 7282 8780 7288 8832
rect 7340 8780 7346 8832
rect 8110 8780 8116 8832
rect 8168 8780 8174 8832
rect 11422 8780 11428 8832
rect 11480 8780 11486 8832
rect 1104 8730 13340 8752
rect 1104 8678 3139 8730
rect 3191 8678 3203 8730
rect 3255 8678 3267 8730
rect 3319 8678 3331 8730
rect 3383 8678 3395 8730
rect 3447 8678 6198 8730
rect 6250 8678 6262 8730
rect 6314 8678 6326 8730
rect 6378 8678 6390 8730
rect 6442 8678 6454 8730
rect 6506 8678 9257 8730
rect 9309 8678 9321 8730
rect 9373 8678 9385 8730
rect 9437 8678 9449 8730
rect 9501 8678 9513 8730
rect 9565 8678 12316 8730
rect 12368 8678 12380 8730
rect 12432 8678 12444 8730
rect 12496 8678 12508 8730
rect 12560 8678 12572 8730
rect 12624 8678 13340 8730
rect 1104 8656 13340 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 2038 8616 2044 8628
rect 1544 8588 2044 8616
rect 1544 8576 1550 8588
rect 2038 8576 2044 8588
rect 2096 8616 2102 8628
rect 2096 8588 2774 8616
rect 2096 8576 2102 8588
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8548 2467 8551
rect 2746 8548 2774 8588
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3016 8588 3249 8616
rect 3016 8576 3022 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3329 8619 3387 8625
rect 3329 8585 3341 8619
rect 3375 8616 3387 8619
rect 3602 8616 3608 8628
rect 3375 8588 3608 8616
rect 3375 8585 3387 8588
rect 3329 8579 3387 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 7282 8616 7288 8628
rect 6135 8588 7288 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 10502 8576 10508 8628
rect 10560 8576 10566 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 3513 8551 3571 8557
rect 2455 8520 2636 8548
rect 2746 8520 3004 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2332 8344 2360 8443
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2608 8489 2636 8520
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2774 8440 2780 8492
rect 2832 8440 2838 8492
rect 2866 8440 2872 8492
rect 2924 8440 2930 8492
rect 2976 8489 3004 8520
rect 3513 8517 3525 8551
rect 3559 8548 3571 8551
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3559 8520 3985 8548
rect 3559 8517 3571 8520
rect 3513 8511 3571 8517
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 4356 8548 4384 8576
rect 4356 8520 4476 8548
rect 3973 8511 4031 8517
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3326 8480 3332 8492
rect 3007 8452 3332 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 3936 8452 4169 8480
rect 3936 8440 3942 8452
rect 4157 8449 4169 8452
rect 4203 8480 4215 8483
rect 4246 8480 4252 8492
rect 4203 8452 4252 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4448 8489 4476 8520
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 6052 8520 6377 8548
rect 6052 8508 6058 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 3050 8412 3056 8424
rect 2746 8384 3056 8412
rect 2746 8344 2774 8384
rect 3050 8372 3056 8384
rect 3108 8412 3114 8424
rect 4448 8412 4476 8443
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5684 8452 5917 8480
rect 5684 8440 5690 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 8294 8480 8300 8492
rect 6227 8452 8300 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 3108 8384 4476 8412
rect 5920 8412 5948 8443
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 10520 8412 10548 8576
rect 12176 8548 12204 8576
rect 12345 8551 12403 8557
rect 12345 8548 12357 8551
rect 12176 8520 12357 8548
rect 12345 8517 12357 8520
rect 12391 8517 12403 8551
rect 12345 8511 12403 8517
rect 12066 8440 12072 8492
rect 12124 8440 12130 8492
rect 5920 8384 10548 8412
rect 3108 8372 3114 8384
rect 12894 8372 12900 8424
rect 12952 8372 12958 8424
rect 2332 8316 2774 8344
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4062 8344 4068 8356
rect 3927 8316 4068 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 12161 8347 12219 8353
rect 12161 8313 12173 8347
rect 12207 8344 12219 8347
rect 12207 8316 12480 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 12452 8288 12480 8316
rect 2222 8236 2228 8288
rect 2280 8276 2286 8288
rect 2774 8276 2780 8288
rect 2280 8248 2780 8276
rect 2280 8236 2286 8248
rect 2774 8236 2780 8248
rect 2832 8276 2838 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 2832 8248 3525 8276
rect 2832 8236 2838 8248
rect 3513 8245 3525 8248
rect 3559 8276 3571 8279
rect 4614 8276 4620 8288
rect 3559 8248 4620 8276
rect 3559 8245 3571 8248
rect 3513 8239 3571 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 7650 8236 7656 8288
rect 7708 8236 7714 8288
rect 12434 8236 12440 8288
rect 12492 8236 12498 8288
rect 1104 8186 13340 8208
rect 1104 8134 2479 8186
rect 2531 8134 2543 8186
rect 2595 8134 2607 8186
rect 2659 8134 2671 8186
rect 2723 8134 2735 8186
rect 2787 8134 5538 8186
rect 5590 8134 5602 8186
rect 5654 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 8597 8186
rect 8649 8134 8661 8186
rect 8713 8134 8725 8186
rect 8777 8134 8789 8186
rect 8841 8134 8853 8186
rect 8905 8134 11656 8186
rect 11708 8134 11720 8186
rect 11772 8134 11784 8186
rect 11836 8134 11848 8186
rect 11900 8134 11912 8186
rect 11964 8134 13340 8186
rect 1104 8112 13340 8134
rect 2222 8032 2228 8084
rect 2280 8032 2286 8084
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 2866 8072 2872 8084
rect 2639 8044 2872 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 2240 7945 2268 8032
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 2406 7828 2412 7880
rect 2464 7828 2470 7880
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2608 7868 2636 8035
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3050 8032 3056 8084
rect 3108 8032 3114 8084
rect 4338 8032 4344 8084
rect 4396 8032 4402 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5132 8044 5549 8072
rect 5132 8032 5138 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 12894 8032 12900 8084
rect 12952 8032 12958 8084
rect 4356 7936 4384 8032
rect 2792 7908 4384 7936
rect 2547 7840 2636 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 2792 7877 2820 7908
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 9180 7908 9321 7936
rect 9180 7896 9186 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 11422 7896 11428 7948
rect 11480 7896 11486 7948
rect 2777 7871 2835 7877
rect 2777 7868 2789 7871
rect 2740 7840 2789 7868
rect 2740 7828 2746 7840
rect 2777 7837 2789 7840
rect 2823 7868 2835 7871
rect 2823 7840 2877 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 3016 7840 3249 7868
rect 3016 7828 3022 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7650 7868 7656 7880
rect 7064 7840 7656 7868
rect 7064 7828 7070 7840
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8478 7868 8484 7880
rect 8251 7840 8484 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9950 7868 9956 7880
rect 9723 7840 9956 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 11146 7828 11152 7880
rect 11204 7828 11210 7880
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2700 7800 2728 7828
rect 8128 7800 8156 7828
rect 2372 7772 2728 7800
rect 6564 7772 8156 7800
rect 2372 7760 2378 7772
rect 6564 7744 6592 7772
rect 8938 7760 8944 7812
rect 8996 7760 9002 7812
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 10134 7800 10140 7812
rect 9171 7772 10140 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 12434 7760 12440 7812
rect 12492 7760 12498 7812
rect 2222 7692 2228 7744
rect 2280 7692 2286 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 8018 7692 8024 7744
rect 8076 7692 8082 7744
rect 8386 7692 8392 7744
rect 8444 7692 8450 7744
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9582 7732 9588 7744
rect 9539 7704 9588 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 1104 7642 13340 7664
rect 1104 7590 3139 7642
rect 3191 7590 3203 7642
rect 3255 7590 3267 7642
rect 3319 7590 3331 7642
rect 3383 7590 3395 7642
rect 3447 7590 6198 7642
rect 6250 7590 6262 7642
rect 6314 7590 6326 7642
rect 6378 7590 6390 7642
rect 6442 7590 6454 7642
rect 6506 7590 9257 7642
rect 9309 7590 9321 7642
rect 9373 7590 9385 7642
rect 9437 7590 9449 7642
rect 9501 7590 9513 7642
rect 9565 7590 12316 7642
rect 12368 7590 12380 7642
rect 12432 7590 12444 7642
rect 12496 7590 12508 7642
rect 12560 7590 12572 7642
rect 12624 7590 13340 7642
rect 1104 7568 13340 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2464 7500 2697 7528
rect 2464 7488 2470 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 2685 7491 2743 7497
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 5951 7500 6224 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 5767 7432 5948 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 5920 7404 5948 7432
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2682 7392 2688 7404
rect 2639 7364 2688 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2958 7392 2964 7404
rect 2823 7364 2964 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6196 7401 6224 7500
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 9232 7500 11192 7528
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 8404 7460 8432 7488
rect 8757 7463 8815 7469
rect 8757 7460 8769 7463
rect 8404 7432 8769 7460
rect 8757 7429 8769 7432
rect 8803 7429 8815 7463
rect 8757 7423 8815 7429
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9232 7401 9260 7500
rect 11164 7472 11192 7500
rect 9493 7463 9551 7469
rect 9493 7429 9505 7463
rect 9539 7460 9551 7463
rect 9582 7460 9588 7472
rect 9539 7432 9588 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 11146 7420 11152 7472
rect 11204 7420 11210 7472
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 9088 7364 9229 7392
rect 9088 7352 9094 7364
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 11241 7395 11299 7401
rect 9217 7355 9275 7361
rect 3528 7324 3556 7352
rect 6564 7324 6592 7352
rect 3528 7296 6592 7324
rect 10612 7324 10640 7378
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 12066 7392 12072 7404
rect 11287 7364 12072 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10612 7296 11161 7324
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11256 7324 11284 7355
rect 12066 7352 12072 7364
rect 12124 7392 12130 7404
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 12124 7364 12173 7392
rect 12124 7352 12130 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 11422 7324 11428 7336
rect 11256 7296 11428 7324
rect 11149 7287 11207 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 4982 7216 4988 7268
rect 5040 7256 5046 7268
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 5040 7228 5365 7256
rect 5040 7216 5046 7228
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 5920 7228 6592 7256
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 4672 7160 5733 7188
rect 4672 7148 4678 7160
rect 5721 7157 5733 7160
rect 5767 7188 5779 7191
rect 5920 7188 5948 7228
rect 6564 7200 6592 7228
rect 5767 7160 5948 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 5994 7148 6000 7200
rect 6052 7148 6058 7200
rect 6546 7148 6552 7200
rect 6604 7148 6610 7200
rect 6641 7191 6699 7197
rect 6641 7157 6653 7191
rect 6687 7188 6699 7191
rect 6914 7188 6920 7200
rect 6687 7160 6920 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7282 7148 7288 7200
rect 7340 7148 7346 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10192 7160 10977 7188
rect 10192 7148 10198 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12434 7188 12440 7200
rect 12299 7160 12440 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 1104 7098 13340 7120
rect 1104 7046 2479 7098
rect 2531 7046 2543 7098
rect 2595 7046 2607 7098
rect 2659 7046 2671 7098
rect 2723 7046 2735 7098
rect 2787 7046 5538 7098
rect 5590 7046 5602 7098
rect 5654 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 8597 7098
rect 8649 7046 8661 7098
rect 8713 7046 8725 7098
rect 8777 7046 8789 7098
rect 8841 7046 8853 7098
rect 8905 7046 11656 7098
rect 11708 7046 11720 7098
rect 11772 7046 11784 7098
rect 11836 7046 11848 7098
rect 11900 7046 11912 7098
rect 11964 7046 13340 7098
rect 1104 7024 13340 7046
rect 1660 6987 1718 6993
rect 1660 6953 1672 6987
rect 1706 6984 1718 6987
rect 2222 6984 2228 6996
rect 1706 6956 2228 6984
rect 1706 6953 1718 6956
rect 1660 6947 1718 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 5800 6987 5858 6993
rect 5800 6953 5812 6987
rect 5846 6984 5858 6987
rect 5994 6984 6000 6996
rect 5846 6956 6000 6984
rect 5846 6953 5858 6956
rect 5800 6947 5858 6953
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 6604 6956 8401 6984
rect 6604 6944 6610 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 8389 6947 8447 6953
rect 8404 6916 8432 6947
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 8573 6987 8631 6993
rect 8573 6984 8585 6987
rect 8536 6956 8585 6984
rect 8536 6944 8542 6956
rect 8573 6953 8585 6956
rect 8619 6953 8631 6987
rect 9309 6987 9367 6993
rect 9309 6984 9321 6987
rect 8573 6947 8631 6953
rect 8680 6956 9321 6984
rect 8680 6916 8708 6956
rect 9309 6953 9321 6956
rect 9355 6953 9367 6987
rect 9309 6947 9367 6953
rect 8404 6888 8708 6916
rect 9125 6919 9183 6925
rect 9125 6885 9137 6919
rect 9171 6885 9183 6919
rect 9324 6916 9352 6947
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9953 6987 10011 6993
rect 9953 6984 9965 6987
rect 9640 6956 9965 6984
rect 9640 6944 9646 6956
rect 9953 6953 9965 6956
rect 9999 6953 10011 6987
rect 9953 6947 10011 6953
rect 10597 6987 10655 6993
rect 10597 6953 10609 6987
rect 10643 6984 10655 6987
rect 10962 6984 10968 6996
rect 10643 6956 10968 6984
rect 10643 6953 10655 6956
rect 10597 6947 10655 6953
rect 10612 6916 10640 6947
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 9324 6888 10640 6916
rect 9125 6879 9183 6885
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4212 6820 5028 6848
rect 4212 6808 4218 6820
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 3108 6752 3433 6780
rect 3108 6740 3114 6752
rect 3421 6749 3433 6752
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4890 6740 4896 6792
rect 4948 6740 4954 6792
rect 5000 6780 5028 6820
rect 5074 6808 5080 6860
rect 5132 6848 5138 6860
rect 5442 6848 5448 6860
rect 5132 6820 5448 6848
rect 5132 6808 5138 6820
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5500 6820 5549 6848
rect 5500 6808 5506 6820
rect 5537 6817 5549 6820
rect 5583 6848 5595 6851
rect 9140 6848 9168 6879
rect 9950 6848 9956 6860
rect 5583 6820 9076 6848
rect 9140 6820 9956 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 9048 6792 9076 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 10468 6820 12909 6848
rect 10468 6808 10474 6820
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 5166 6780 5172 6792
rect 5000 6752 5172 6780
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7340 6752 7573 6780
rect 7340 6740 7346 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7975 6752 8033 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8021 6749 8033 6752
rect 8067 6780 8079 6783
rect 8938 6780 8944 6792
rect 8067 6752 8944 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 2898 6684 3341 6712
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 3329 6675 3387 6681
rect 3694 6672 3700 6724
rect 3752 6712 3758 6724
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 3752 6684 4169 6712
rect 3752 6672 3758 6684
rect 4157 6681 4169 6684
rect 4203 6681 4215 6715
rect 4157 6675 4215 6681
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4341 6715 4399 6721
rect 4341 6712 4353 6715
rect 4304 6684 4353 6712
rect 4304 6672 4310 6684
rect 4341 6681 4353 6684
rect 4387 6681 4399 6715
rect 4341 6675 4399 6681
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 5077 6715 5135 6721
rect 5077 6712 5089 6715
rect 4488 6684 5089 6712
rect 4488 6672 4494 6684
rect 5077 6681 5089 6684
rect 5123 6681 5135 6715
rect 5077 6675 5135 6681
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5350 6712 5356 6724
rect 5307 6684 5356 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 5902 6712 5908 6724
rect 5491 6684 5908 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7760 6712 7788 6743
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9030 6740 9036 6792
rect 9088 6740 9094 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9677 6783 9735 6789
rect 9180 6752 9352 6780
rect 9180 6740 9186 6752
rect 9324 6721 9352 6752
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 7248 6684 7788 6712
rect 9309 6715 9367 6721
rect 7248 6672 7254 6684
rect 9309 6681 9321 6715
rect 9355 6681 9367 6715
rect 9309 6675 9367 6681
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 3016 6616 3157 6644
rect 3016 6604 3022 6616
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3145 6607 3203 6613
rect 4522 6604 4528 6656
rect 4580 6604 4586 6656
rect 4706 6604 4712 6656
rect 4764 6604 4770 6656
rect 5368 6644 5396 6672
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 5368 6616 7297 6644
rect 7285 6613 7297 6616
rect 7331 6644 7343 6647
rect 7374 6644 7380 6656
rect 7331 6616 7380 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 9692 6644 9720 6743
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 9916 6752 10241 6780
rect 9916 6740 9922 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10873 6783 10931 6789
rect 10873 6780 10885 6783
rect 10229 6743 10287 6749
rect 10796 6752 10885 6780
rect 9784 6712 9812 6740
rect 9784 6684 9904 6712
rect 9766 6644 9772 6656
rect 9692 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 9876 6644 9904 6684
rect 10134 6672 10140 6724
rect 10192 6672 10198 6724
rect 9937 6647 9995 6653
rect 9937 6644 9949 6647
rect 9876 6616 9949 6644
rect 9937 6613 9949 6616
rect 9983 6613 9995 6647
rect 9937 6607 9995 6613
rect 10594 6604 10600 6656
rect 10652 6604 10658 6656
rect 10796 6653 10824 6752
rect 10873 6749 10885 6752
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11146 6740 11152 6792
rect 11204 6740 11210 6792
rect 11425 6715 11483 6721
rect 11425 6712 11437 6715
rect 11072 6684 11437 6712
rect 11072 6653 11100 6684
rect 11425 6681 11437 6684
rect 11471 6681 11483 6715
rect 11425 6675 11483 6681
rect 12434 6672 12440 6724
rect 12492 6672 12498 6724
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6613 10839 6647
rect 10781 6607 10839 6613
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6613 11115 6647
rect 11057 6607 11115 6613
rect 1104 6554 13340 6576
rect 1104 6502 3139 6554
rect 3191 6502 3203 6554
rect 3255 6502 3267 6554
rect 3319 6502 3331 6554
rect 3383 6502 3395 6554
rect 3447 6502 6198 6554
rect 6250 6502 6262 6554
rect 6314 6502 6326 6554
rect 6378 6502 6390 6554
rect 6442 6502 6454 6554
rect 6506 6502 9257 6554
rect 9309 6502 9321 6554
rect 9373 6502 9385 6554
rect 9437 6502 9449 6554
rect 9501 6502 9513 6554
rect 9565 6502 12316 6554
rect 12368 6502 12380 6554
rect 12432 6502 12444 6554
rect 12496 6502 12508 6554
rect 12560 6502 12572 6554
rect 12624 6502 13340 6554
rect 1104 6480 13340 6502
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 4430 6440 4436 6452
rect 3927 6412 4436 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 7190 6440 7196 6452
rect 5040 6412 7196 6440
rect 5040 6400 5046 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8444 6412 8585 6440
rect 8444 6400 8450 6412
rect 8573 6409 8585 6412
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 9674 6440 9680 6452
rect 8720 6412 9680 6440
rect 8720 6400 8726 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 9824 6412 9996 6440
rect 9824 6400 9830 6412
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 1452 6344 3464 6372
rect 1452 6332 1458 6344
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 2869 6307 2927 6313
rect 2639 6276 2774 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2314 6196 2320 6248
rect 2372 6196 2378 6248
rect 2746 6236 2774 6276
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 3142 6304 3148 6316
rect 2915 6276 3148 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3050 6236 3056 6248
rect 2746 6208 3056 6236
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 2332 6168 2360 6196
rect 3160 6168 3188 6264
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6205 3387 6239
rect 3436 6236 3464 6344
rect 4019 6341 4077 6347
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6304 3571 6307
rect 4019 6307 4031 6341
rect 4065 6338 4077 6341
rect 4065 6307 4092 6338
rect 4246 6332 4252 6384
rect 4304 6332 4310 6384
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6372 4675 6375
rect 4724 6372 4752 6400
rect 5902 6372 5908 6384
rect 4663 6344 4752 6372
rect 5842 6344 5908 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 4019 6304 4092 6307
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 3559 6276 4092 6304
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 4064 6248 4092 6276
rect 4172 6276 4353 6304
rect 3436 6208 3556 6236
rect 3329 6199 3387 6205
rect 2332 6140 3188 6168
rect 3344 6168 3372 6199
rect 3528 6168 3556 6208
rect 3694 6196 3700 6248
rect 3752 6196 3758 6248
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 4172 6168 4200 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 7208 6304 7236 6400
rect 7282 6332 7288 6384
rect 7340 6372 7346 6384
rect 7340 6344 8616 6372
rect 7340 6332 7346 6344
rect 8404 6313 8432 6344
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 7208 6276 8217 6304
rect 4341 6267 4399 6273
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8588 6304 8616 6344
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 9493 6375 9551 6381
rect 9493 6372 9505 6375
rect 9180 6344 9505 6372
rect 9180 6332 9186 6344
rect 9493 6341 9505 6344
rect 9539 6372 9551 6375
rect 9539 6344 9812 6372
rect 9539 6341 9551 6344
rect 9493 6335 9551 6341
rect 9582 6304 9588 6316
rect 8588 6276 9588 6304
rect 8389 6267 8447 6273
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 5258 6236 5264 6248
rect 4304 6208 5264 6236
rect 4304 6196 4310 6208
rect 5258 6196 5264 6208
rect 5316 6236 5322 6248
rect 6089 6239 6147 6245
rect 6089 6236 6101 6239
rect 5316 6208 6101 6236
rect 5316 6196 5322 6208
rect 6089 6205 6101 6208
rect 6135 6205 6147 6239
rect 8220 6236 8248 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9784 6304 9812 6344
rect 9858 6332 9864 6384
rect 9916 6332 9922 6384
rect 9968 6381 9996 6412
rect 10042 6400 10048 6452
rect 10100 6400 10106 6452
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10594 6440 10600 6452
rect 10367 6412 10600 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 9953 6375 10011 6381
rect 9953 6341 9965 6375
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 10060 6304 10088 6400
rect 10137 6375 10195 6381
rect 10137 6341 10149 6375
rect 10183 6372 10195 6375
rect 10410 6372 10416 6384
rect 10183 6344 10416 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 9784 6276 10088 6304
rect 8662 6236 8668 6248
rect 8220 6208 8668 6236
rect 6089 6199 6147 6205
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6236 9367 6239
rect 9766 6236 9772 6248
rect 9355 6208 9772 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9766 6196 9772 6208
rect 9824 6236 9830 6248
rect 10152 6236 10180 6335
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12032 6276 12725 6304
rect 12032 6264 12038 6276
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 9824 6208 10180 6236
rect 9824 6196 9830 6208
rect 12986 6196 12992 6248
rect 13044 6196 13050 6248
rect 3344 6140 3464 6168
rect 3528 6140 4200 6168
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2188 6072 2421 6100
rect 2188 6060 2194 6072
rect 2409 6069 2421 6072
rect 2455 6069 2467 6103
rect 2409 6063 2467 6069
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2866 6100 2872 6112
rect 2823 6072 2872 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3436 6100 3464 6140
rect 3970 6100 3976 6112
rect 3436 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 4028 6072 4077 6100
rect 4028 6060 4034 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4172 6100 4200 6140
rect 5074 6100 5080 6112
rect 4172 6072 5080 6100
rect 4065 6063 4123 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 1104 6010 13340 6032
rect 1104 5958 2479 6010
rect 2531 5958 2543 6010
rect 2595 5958 2607 6010
rect 2659 5958 2671 6010
rect 2723 5958 2735 6010
rect 2787 5958 5538 6010
rect 5590 5958 5602 6010
rect 5654 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 8597 6010
rect 8649 5958 8661 6010
rect 8713 5958 8725 6010
rect 8777 5958 8789 6010
rect 8841 5958 8853 6010
rect 8905 5958 11656 6010
rect 11708 5958 11720 6010
rect 11772 5958 11784 6010
rect 11836 5958 11848 6010
rect 11900 5958 11912 6010
rect 11964 5958 13340 6010
rect 1104 5936 13340 5958
rect 1394 5856 1400 5908
rect 1452 5856 1458 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 4430 5856 4436 5908
rect 4488 5856 4494 5908
rect 4522 5856 4528 5908
rect 4580 5856 4586 5908
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 5224 5868 6469 5896
rect 5224 5856 5230 5868
rect 6457 5865 6469 5868
rect 6503 5896 6515 5899
rect 6914 5896 6920 5908
rect 6503 5868 6920 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 1412 5760 1440 5856
rect 3973 5831 4031 5837
rect 3973 5797 3985 5831
rect 4019 5828 4031 5831
rect 4448 5828 4476 5856
rect 4019 5800 4476 5828
rect 4019 5797 4031 5800
rect 3973 5791 4031 5797
rect 1489 5763 1547 5769
rect 1489 5760 1501 5763
rect 1412 5732 1501 5760
rect 1489 5729 1501 5732
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 2130 5760 2136 5772
rect 1811 5732 2136 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2866 5652 2872 5704
rect 2924 5652 2930 5704
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 4540 5624 4568 5856
rect 4387 5596 4568 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3970 5556 3976 5568
rect 3283 5528 3976 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4525 5559 4583 5565
rect 4525 5525 4537 5559
rect 4571 5556 4583 5559
rect 4908 5556 4936 5856
rect 8754 5828 8760 5840
rect 8128 5800 8760 5828
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8128 5760 8156 5800
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 7975 5732 8156 5760
rect 8205 5763 8263 5769
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 9030 5760 9036 5772
rect 8251 5732 9036 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 8220 5664 8309 5692
rect 8220 5636 8248 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 6365 5627 6423 5633
rect 6365 5593 6377 5627
rect 6411 5624 6423 5627
rect 6411 5596 6684 5624
rect 7498 5596 7604 5624
rect 6411 5593 6423 5596
rect 6365 5587 6423 5593
rect 4571 5528 4936 5556
rect 6656 5556 6684 5596
rect 7006 5556 7012 5568
rect 6656 5528 7012 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7576 5556 7604 5596
rect 8202 5584 8208 5636
rect 8260 5584 8266 5636
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 8404 5556 8432 5587
rect 7576 5528 8432 5556
rect 1104 5466 13340 5488
rect 1104 5414 3139 5466
rect 3191 5414 3203 5466
rect 3255 5414 3267 5466
rect 3319 5414 3331 5466
rect 3383 5414 3395 5466
rect 3447 5414 6198 5466
rect 6250 5414 6262 5466
rect 6314 5414 6326 5466
rect 6378 5414 6390 5466
rect 6442 5414 6454 5466
rect 6506 5414 9257 5466
rect 9309 5414 9321 5466
rect 9373 5414 9385 5466
rect 9437 5414 9449 5466
rect 9501 5414 9513 5466
rect 9565 5414 12316 5466
rect 12368 5414 12380 5466
rect 12432 5414 12444 5466
rect 12496 5414 12508 5466
rect 12560 5414 12572 5466
rect 12624 5414 13340 5466
rect 1104 5392 13340 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 3050 5352 3056 5364
rect 2823 5324 3056 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 4982 5312 4988 5364
rect 5040 5312 5046 5364
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5316 5324 5365 5352
rect 5316 5312 5322 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5902 5352 5908 5364
rect 5767 5324 5908 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 8754 5312 8760 5364
rect 8812 5312 8818 5364
rect 9122 5312 9128 5364
rect 9180 5312 9186 5364
rect 9766 5312 9772 5364
rect 9824 5312 9830 5364
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 11333 5355 11391 5361
rect 10459 5324 11008 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 2314 5244 2320 5296
rect 2372 5284 2378 5296
rect 2409 5287 2467 5293
rect 2409 5284 2421 5287
rect 2372 5256 2421 5284
rect 2372 5244 2378 5256
rect 2409 5253 2421 5256
rect 2455 5253 2467 5287
rect 2409 5247 2467 5253
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 3007 5256 3801 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 3789 5253 3801 5256
rect 3835 5253 3847 5287
rect 3789 5247 3847 5253
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2148 5024 2176 5179
rect 2424 5148 2452 5247
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 4157 5287 4215 5293
rect 4157 5284 4169 5287
rect 4120 5256 4169 5284
rect 4120 5244 4126 5256
rect 4157 5253 4169 5256
rect 4203 5284 4215 5287
rect 5169 5287 5227 5293
rect 5169 5284 5181 5287
rect 4203 5256 5181 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 5169 5253 5181 5256
rect 5215 5253 5227 5287
rect 5169 5247 5227 5253
rect 5534 5244 5540 5296
rect 5592 5244 5598 5296
rect 8294 5293 8300 5296
rect 8271 5287 8300 5293
rect 8271 5253 8283 5287
rect 8271 5247 8300 5253
rect 8294 5244 8300 5247
rect 8352 5244 8358 5296
rect 9140 5284 9168 5312
rect 9140 5256 9352 5284
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3694 5216 3700 5228
rect 3375 5188 3700 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4028 5188 5273 5216
rect 4028 5176 4034 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5828 5148 5856 5179
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 6972 5188 7389 5216
rect 6972 5176 6978 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 2424 5120 5856 5148
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 8067 5120 8125 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8404 5148 8432 5179
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 9214 5216 9220 5228
rect 8619 5188 9220 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9324 5225 9352 5256
rect 9784 5225 9812 5312
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5185 9827 5219
rect 9876 5216 9904 5312
rect 10505 5287 10563 5293
rect 10505 5284 10517 5287
rect 10244 5256 10517 5284
rect 10244 5225 10272 5256
rect 10505 5253 10517 5256
rect 10551 5253 10563 5287
rect 10505 5247 10563 5253
rect 10686 5244 10692 5296
rect 10744 5244 10750 5296
rect 10980 5293 11008 5324
rect 11333 5321 11345 5355
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 10965 5287 11023 5293
rect 10965 5253 10977 5287
rect 11011 5253 11023 5287
rect 10965 5247 11023 5253
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9876 5188 10241 5216
rect 9769 5179 9827 5185
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 10704 5216 10732 5244
rect 10459 5188 10732 5216
rect 10980 5216 11008 5247
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11165 5287 11223 5293
rect 11165 5284 11177 5287
rect 11112 5256 11177 5284
rect 11112 5244 11118 5256
rect 11165 5253 11177 5256
rect 11211 5253 11223 5287
rect 11165 5247 11223 5253
rect 11348 5216 11376 5315
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 10980 5188 11284 5216
rect 11348 5188 11713 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 9858 5148 9864 5160
rect 8352 5120 9864 5148
rect 8352 5108 8358 5120
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 11256 5024 11284 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5185 12219 5219
rect 12161 5179 12219 5185
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 12176 5148 12204 5179
rect 11480 5120 12204 5148
rect 11480 5108 11486 5120
rect 2130 4972 2136 5024
rect 2188 4972 2194 5024
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 4338 5012 4344 5024
rect 3007 4984 4344 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 9217 5015 9275 5021
rect 9217 5012 9229 5015
rect 8260 4984 9229 5012
rect 8260 4972 8266 4984
rect 9217 4981 9229 4984
rect 9263 4981 9275 5015
rect 9217 4975 9275 4981
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 9766 5012 9772 5024
rect 9723 4984 9772 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10873 5015 10931 5021
rect 10873 4981 10885 5015
rect 10919 5012 10931 5015
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 10919 4984 11161 5012
rect 10919 4981 10931 4984
rect 10873 4975 10931 4981
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 11238 4972 11244 5024
rect 11296 4972 11302 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 12216 4984 12265 5012
rect 12216 4972 12222 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 1104 4922 13340 4944
rect 1104 4870 2479 4922
rect 2531 4870 2543 4922
rect 2595 4870 2607 4922
rect 2659 4870 2671 4922
rect 2723 4870 2735 4922
rect 2787 4870 5538 4922
rect 5590 4870 5602 4922
rect 5654 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 8597 4922
rect 8649 4870 8661 4922
rect 8713 4870 8725 4922
rect 8777 4870 8789 4922
rect 8841 4870 8853 4922
rect 8905 4870 11656 4922
rect 11708 4870 11720 4922
rect 11772 4870 11784 4922
rect 11836 4870 11848 4922
rect 11900 4870 11912 4922
rect 11964 4870 13340 4922
rect 1104 4848 13340 4870
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 9272 4780 10701 4808
rect 9272 4768 9278 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 11422 4808 11428 4820
rect 10689 4771 10747 4777
rect 11256 4780 11428 4808
rect 11256 4740 11284 4780
rect 11422 4768 11428 4780
rect 11480 4808 11486 4820
rect 12802 4808 12808 4820
rect 11480 4780 12808 4808
rect 11480 4768 11486 4780
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 4816 4712 11284 4740
rect 4816 4684 4844 4712
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4672 3019 4675
rect 4798 4672 4804 4684
rect 3007 4644 4804 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11514 4672 11520 4684
rect 11471 4644 11520 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 2130 4468 2136 4480
rect 1627 4440 2136 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 2130 4428 2136 4440
rect 2188 4468 2194 4480
rect 2700 4468 2728 4567
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 10919 4576 11100 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 10704 4536 10732 4564
rect 10962 4536 10968 4548
rect 10704 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11072 4480 11100 4576
rect 11146 4564 11152 4616
rect 11204 4564 11210 4616
rect 12158 4496 12164 4548
rect 12216 4496 12222 4548
rect 2188 4440 2728 4468
rect 2188 4428 2194 4440
rect 11054 4428 11060 4480
rect 11112 4428 11118 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 11388 4440 12909 4468
rect 11388 4428 11394 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 1104 4378 13340 4400
rect 1104 4326 3139 4378
rect 3191 4326 3203 4378
rect 3255 4326 3267 4378
rect 3319 4326 3331 4378
rect 3383 4326 3395 4378
rect 3447 4326 6198 4378
rect 6250 4326 6262 4378
rect 6314 4326 6326 4378
rect 6378 4326 6390 4378
rect 6442 4326 6454 4378
rect 6506 4326 9257 4378
rect 9309 4326 9321 4378
rect 9373 4326 9385 4378
rect 9437 4326 9449 4378
rect 9501 4326 9513 4378
rect 9565 4326 12316 4378
rect 12368 4326 12380 4378
rect 12432 4326 12444 4378
rect 12496 4326 12508 4378
rect 12560 4326 12572 4378
rect 12624 4326 13340 4378
rect 1104 4304 13340 4326
rect 2792 4236 3188 4264
rect 2792 4128 2820 4236
rect 2056 4100 2820 4128
rect 2869 4131 2927 4137
rect 2056 4072 2084 4100
rect 2869 4097 2881 4131
rect 2915 4097 2927 4131
rect 3160 4128 3188 4236
rect 3326 4224 3332 4276
rect 3384 4224 3390 4276
rect 4154 4224 4160 4276
rect 4212 4224 4218 4276
rect 4448 4236 6224 4264
rect 4338 4128 4344 4140
rect 3160 4100 4344 4128
rect 2869 4091 2927 4097
rect 2038 4020 2044 4072
rect 2096 4020 2102 4072
rect 2222 4020 2228 4072
rect 2280 4060 2286 4072
rect 2682 4060 2688 4072
rect 2280 4032 2688 4060
rect 2280 4020 2286 4032
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 2884 4060 2912 4091
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 3694 4060 3700 4072
rect 2884 4032 3700 4060
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 4448 4060 4476 4236
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5994 4196 6000 4208
rect 5675 4168 6000 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4571 4100 4660 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 3804 4032 4476 4060
rect 4632 4060 4660 4100
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5123 4100 5733 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 6196 4128 6224 4236
rect 7190 4224 7196 4276
rect 7248 4224 7254 4276
rect 7282 4224 7288 4276
rect 7340 4224 7346 4276
rect 10229 4267 10287 4273
rect 7668 4236 9076 4264
rect 7208 4137 7236 4224
rect 7300 4196 7328 4224
rect 7668 4205 7696 4236
rect 7653 4199 7711 4205
rect 7653 4196 7665 4199
rect 7300 4168 7665 4196
rect 7653 4165 7665 4168
rect 7699 4165 7711 4199
rect 7653 4159 7711 4165
rect 7944 4168 8524 4196
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6196 4100 6929 4128
rect 5721 4091 5779 4097
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7374 4088 7380 4140
rect 7432 4088 7438 4140
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 5350 4060 5356 4072
rect 4632 4032 5356 4060
rect 2593 3995 2651 4001
rect 2593 3961 2605 3995
rect 2639 3992 2651 3995
rect 3050 3992 3056 4004
rect 2639 3964 3056 3992
rect 2639 3961 2651 3964
rect 2593 3955 2651 3961
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 3804 3992 3832 4032
rect 3660 3964 3832 3992
rect 3660 3952 3666 3964
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 4065 3995 4123 4001
rect 4065 3992 4077 3995
rect 4028 3964 4077 3992
rect 4028 3952 4034 3964
rect 4065 3961 4077 3964
rect 4111 3992 4123 3995
rect 4632 3992 4660 4032
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 5902 4060 5908 4072
rect 5859 4032 5908 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 6086 4060 6092 4072
rect 6043 4032 6092 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6512 4032 6745 4060
rect 6512 4020 6518 4032
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7944 4060 7972 4168
rect 8018 4088 8024 4140
rect 8076 4088 8082 4140
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 8168 4100 8217 4128
rect 8168 4088 8174 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 6880 4032 7972 4060
rect 8312 4060 8340 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8496 4128 8524 4168
rect 8772 4168 8984 4196
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8496 4100 8677 4128
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8772 4060 8800 4168
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 8312 4032 8800 4060
rect 6880 4020 6886 4032
rect 4111 3964 4660 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 5258 3952 5264 4004
rect 5316 3952 5322 4004
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 7009 3995 7067 4001
rect 7009 3992 7021 3995
rect 5500 3964 7021 3992
rect 5500 3952 5506 3964
rect 7009 3961 7021 3964
rect 7055 3961 7067 3995
rect 7009 3955 7067 3961
rect 7098 3952 7104 4004
rect 7156 3952 7162 4004
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 7929 3995 7987 4001
rect 7248 3964 7880 3992
rect 7248 3952 7254 3964
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2866 3924 2872 3936
rect 2731 3896 2872 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 3878 3924 3884 3936
rect 3191 3896 3884 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 5074 3924 5080 3936
rect 4663 3896 5080 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5166 3884 5172 3936
rect 5224 3884 5230 3936
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 6638 3924 6644 3936
rect 5951 3896 6644 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7558 3924 7564 3936
rect 6972 3896 7564 3924
rect 6972 3884 6978 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7852 3924 7880 3964
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8864 3992 8892 4091
rect 8956 4060 8984 4168
rect 9048 4128 9076 4236
rect 10229 4233 10241 4267
rect 10275 4264 10287 4267
rect 10870 4264 10876 4276
rect 10275 4236 10876 4264
rect 10275 4233 10287 4236
rect 10229 4227 10287 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 11330 4264 11336 4276
rect 11020 4236 11336 4264
rect 11020 4224 11026 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11149 4199 11207 4205
rect 11149 4196 11161 4199
rect 11112 4168 11161 4196
rect 11112 4156 11118 4168
rect 11149 4165 11161 4168
rect 11195 4196 11207 4199
rect 11195 4168 12940 4196
rect 11195 4165 11207 4168
rect 11149 4159 11207 4165
rect 12912 4140 12940 4168
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9048 4100 9413 4128
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 9766 4088 9772 4140
rect 9824 4088 9830 4140
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10379 4131 10437 4137
rect 10379 4128 10391 4131
rect 9916 4100 10391 4128
rect 9916 4088 9922 4100
rect 10379 4097 10391 4100
rect 10425 4128 10437 4131
rect 10425 4097 10456 4128
rect 10379 4091 10456 4097
rect 9784 4060 9812 4088
rect 8956 4032 9812 4060
rect 10428 4004 10456 4091
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 11747 4100 12357 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12894 4088 12900 4140
rect 12952 4088 12958 4140
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 7975 3964 8892 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 9122 3952 9128 4004
rect 9180 3952 9186 4004
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9272 3964 10364 3992
rect 9272 3952 9278 3964
rect 8386 3924 8392 3936
rect 7852 3896 8392 3924
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8536 3896 8585 3924
rect 8536 3884 8542 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8573 3887 8631 3893
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 8938 3924 8944 3936
rect 8895 3896 8944 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 9088 3896 9321 3924
rect 9088 3884 9094 3896
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 10336 3924 10364 3964
rect 10410 3952 10416 4004
rect 10468 3952 10474 4004
rect 10796 3992 10824 4023
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11296 4032 11621 4060
rect 11296 4020 11302 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 10796 3964 11161 3992
rect 11149 3961 11161 3964
rect 11195 3961 11207 3995
rect 11149 3955 11207 3961
rect 10778 3924 10784 3936
rect 10336 3896 10784 3924
rect 9309 3887 9367 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 12066 3884 12072 3936
rect 12124 3884 12130 3936
rect 1104 3834 13340 3856
rect 1104 3782 2479 3834
rect 2531 3782 2543 3834
rect 2595 3782 2607 3834
rect 2659 3782 2671 3834
rect 2723 3782 2735 3834
rect 2787 3782 5538 3834
rect 5590 3782 5602 3834
rect 5654 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 8597 3834
rect 8649 3782 8661 3834
rect 8713 3782 8725 3834
rect 8777 3782 8789 3834
rect 8841 3782 8853 3834
rect 8905 3782 11656 3834
rect 11708 3782 11720 3834
rect 11772 3782 11784 3834
rect 11836 3782 11848 3834
rect 11900 3782 11912 3834
rect 11964 3782 13340 3834
rect 1104 3760 13340 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 1719 3692 2329 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 2317 3683 2375 3689
rect 2685 3723 2743 3729
rect 2685 3689 2697 3723
rect 2731 3720 2743 3723
rect 2866 3720 2872 3732
rect 2731 3692 2872 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 1949 3655 2007 3661
rect 1949 3621 1961 3655
rect 1995 3652 2007 3655
rect 2222 3652 2228 3664
rect 1995 3624 2228 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3516 1455 3519
rect 1578 3516 1584 3528
rect 1443 3488 1584 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 1578 3476 1584 3488
rect 1636 3516 1642 3528
rect 1964 3516 1992 3615
rect 2222 3612 2228 3624
rect 2280 3612 2286 3664
rect 2038 3544 2044 3596
rect 2096 3544 2102 3596
rect 2332 3584 2360 3683
rect 2866 3680 2872 3692
rect 2924 3720 2930 3732
rect 4525 3723 4583 3729
rect 2924 3692 4200 3720
rect 2924 3680 2930 3692
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3652 2559 3655
rect 2547 3624 3280 3652
rect 2547 3621 2559 3624
rect 2501 3615 2559 3621
rect 2958 3584 2964 3596
rect 2332 3556 2964 3584
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 1636 3488 1992 3516
rect 2056 3516 2084 3544
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2056 3488 2605 3516
rect 1636 3476 1642 3488
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 2961 3451 3019 3457
rect 2961 3448 2973 3451
rect 1872 3420 2973 3448
rect 1872 3389 1900 3420
rect 2961 3417 2973 3420
rect 3007 3417 3019 3451
rect 3252 3448 3280 3624
rect 3326 3612 3332 3664
rect 3384 3612 3390 3664
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 3559 3624 4108 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 3344 3584 3372 3612
rect 4080 3596 4108 3624
rect 3344 3556 3832 3584
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3602 3516 3608 3528
rect 3467 3488 3608 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 3804 3525 3832 3556
rect 4062 3544 4068 3596
rect 4120 3544 4126 3596
rect 4172 3593 4200 3692
rect 4525 3689 4537 3723
rect 4571 3720 4583 3723
rect 4798 3720 4804 3732
rect 4571 3692 4804 3720
rect 4571 3689 4583 3692
rect 4525 3683 4583 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 6822 3720 6828 3732
rect 5583 3692 6828 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3689 7067 3723
rect 7009 3683 7067 3689
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3553 4215 3587
rect 5092 3584 5120 3680
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 6086 3652 6092 3664
rect 5951 3624 6092 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 6914 3652 6920 3664
rect 6288 3624 6920 3652
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 5092 3556 5181 3584
rect 4157 3547 4215 3553
rect 5169 3553 5181 3556
rect 5215 3584 5227 3587
rect 5442 3584 5448 3596
rect 5215 3556 5448 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 5442 3544 5448 3556
rect 5500 3584 5506 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 5500 3556 5733 3584
rect 5500 3544 5506 3556
rect 5721 3553 5733 3556
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 5994 3544 6000 3596
rect 6052 3544 6058 3596
rect 6288 3584 6316 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7024 3652 7052 3683
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7156 3692 7389 3720
rect 7156 3680 7162 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 8018 3680 8024 3732
rect 8076 3720 8082 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8076 3692 8953 3720
rect 8076 3680 8082 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 9214 3720 9220 3732
rect 8941 3683 8999 3689
rect 9140 3692 9220 3720
rect 7024 3624 8616 3652
rect 6104 3556 6316 3584
rect 6365 3587 6423 3593
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 3988 3448 4016 3479
rect 4338 3476 4344 3528
rect 4396 3476 4402 3528
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 3252 3420 4016 3448
rect 2961 3411 3019 3417
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3349 1915 3383
rect 1857 3343 1915 3349
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 2096 3352 2329 3380
rect 2096 3340 2102 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 2866 3340 2872 3392
rect 2924 3340 2930 3392
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 5000 3380 5028 3479
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 6012 3516 6040 3544
rect 6104 3528 6132 3556
rect 6365 3553 6377 3587
rect 6411 3584 6423 3587
rect 6411 3556 6960 3584
rect 6411 3553 6423 3556
rect 6365 3547 6423 3553
rect 5859 3488 6040 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 5368 3448 5396 3479
rect 6086 3476 6092 3528
rect 6144 3476 6150 3528
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3516 6515 3519
rect 6730 3516 6736 3528
rect 6503 3488 6736 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 6197 3448 6225 3479
rect 5368 3420 6225 3448
rect 3375 3352 5028 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6472 3380 6500 3479
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 6932 3516 6960 3556
rect 7098 3544 7104 3596
rect 7156 3544 7162 3596
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7340 3556 7512 3584
rect 7340 3544 7346 3556
rect 6932 3488 7052 3516
rect 6914 3408 6920 3460
rect 6972 3408 6978 3460
rect 7024 3448 7052 3488
rect 7190 3476 7196 3528
rect 7248 3476 7254 3528
rect 7484 3516 7512 3556
rect 7742 3544 7748 3596
rect 7800 3544 7806 3596
rect 7594 3519 7652 3525
rect 7594 3516 7606 3519
rect 7484 3488 7606 3516
rect 7594 3485 7606 3488
rect 7640 3485 7652 3519
rect 7594 3479 7652 3485
rect 7760 3448 7788 3544
rect 7944 3516 7972 3624
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8478 3584 8484 3596
rect 8067 3556 8484 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 8588 3528 8616 3624
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9140 3584 9168 3692
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 10229 3723 10287 3729
rect 9324 3692 9812 3720
rect 9324 3652 9352 3692
rect 9784 3664 9812 3692
rect 10229 3689 10241 3723
rect 10275 3720 10287 3723
rect 10686 3720 10692 3732
rect 10275 3692 10692 3720
rect 10275 3689 10287 3692
rect 10229 3683 10287 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10928 3692 10977 3720
rect 10928 3680 10934 3692
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 10965 3683 11023 3689
rect 12894 3680 12900 3732
rect 12952 3680 12958 3732
rect 8904 3556 9168 3584
rect 8904 3544 8910 3556
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7944 3488 8125 3516
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8202 3476 8208 3528
rect 8260 3476 8266 3528
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8720 3488 8769 3516
rect 8720 3476 8726 3488
rect 8757 3485 8769 3488
rect 8803 3516 8815 3519
rect 9030 3516 9036 3528
rect 8803 3488 9036 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 9140 3525 9168 3556
rect 9232 3624 9352 3652
rect 9232 3525 9260 3624
rect 9398 3612 9404 3664
rect 9456 3612 9462 3664
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 9640 3612 9674 3652
rect 9766 3612 9772 3664
rect 9824 3612 9830 3664
rect 9646 3584 9674 3612
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 9646 3556 10517 3584
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10888 3584 10916 3680
rect 10505 3547 10563 3553
rect 10612 3556 10916 3584
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9475 3519 9533 3525
rect 9475 3516 9487 3519
rect 9364 3488 9487 3516
rect 9364 3476 9370 3488
rect 9475 3485 9487 3488
rect 9521 3485 9533 3519
rect 9475 3479 9533 3485
rect 9582 3476 9588 3528
rect 9640 3476 9646 3528
rect 9674 3476 9680 3528
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 10612 3525 10640 3556
rect 11146 3544 11152 3596
rect 11204 3544 11210 3596
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9824 3488 9965 3516
rect 9824 3476 9830 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 10050 3519 10108 3525
rect 10050 3485 10062 3519
rect 10096 3516 10108 3519
rect 10413 3519 10471 3525
rect 10096 3488 10180 3516
rect 10096 3485 10108 3488
rect 10050 3479 10108 3485
rect 7024 3420 7788 3448
rect 8220 3448 8248 3476
rect 8481 3451 8539 3457
rect 8481 3448 8493 3451
rect 8220 3420 8493 3448
rect 5868 3352 6500 3380
rect 5868 3340 5874 3352
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 7760 3380 7788 3420
rect 8481 3417 8493 3420
rect 8527 3417 8539 3451
rect 8481 3411 8539 3417
rect 7699 3352 7788 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 8202 3340 8208 3392
rect 8260 3340 8266 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8496 3380 8524 3411
rect 8938 3408 8944 3460
rect 8996 3448 9002 3460
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 8996 3420 9873 3448
rect 8996 3408 9002 3420
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 9861 3411 9919 3417
rect 9030 3380 9036 3392
rect 8352 3352 9036 3380
rect 8352 3340 8358 3352
rect 9030 3340 9036 3352
rect 9088 3380 9094 3392
rect 9306 3380 9312 3392
rect 9088 3352 9312 3380
rect 9088 3340 9094 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10152 3380 10180 3488
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10428 3448 10456 3479
rect 10870 3476 10876 3528
rect 10928 3476 10934 3528
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 10980 3448 11008 3476
rect 10428 3420 11008 3448
rect 11425 3451 11483 3457
rect 11425 3417 11437 3451
rect 11471 3417 11483 3451
rect 12710 3448 12716 3460
rect 12650 3420 12716 3448
rect 11425 3411 11483 3417
rect 11054 3380 11060 3392
rect 9456 3352 11060 3380
rect 9456 3340 9462 3352
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 11440 3380 11468 3411
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 12158 3380 12164 3392
rect 11440 3352 12164 3380
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 1104 3290 13340 3312
rect 1104 3238 3139 3290
rect 3191 3238 3203 3290
rect 3255 3238 3267 3290
rect 3319 3238 3331 3290
rect 3383 3238 3395 3290
rect 3447 3238 6198 3290
rect 6250 3238 6262 3290
rect 6314 3238 6326 3290
rect 6378 3238 6390 3290
rect 6442 3238 6454 3290
rect 6506 3238 9257 3290
rect 9309 3238 9321 3290
rect 9373 3238 9385 3290
rect 9437 3238 9449 3290
rect 9501 3238 9513 3290
rect 9565 3238 12316 3290
rect 12368 3238 12380 3290
rect 12432 3238 12444 3290
rect 12496 3238 12508 3290
rect 12560 3238 12572 3290
rect 12624 3238 13340 3290
rect 1104 3216 13340 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2924 3148 2973 3176
rect 2924 3136 2930 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 3050 3136 3056 3188
rect 3108 3136 3114 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3878 3176 3884 3188
rect 3384 3148 3884 3176
rect 3384 3136 3390 3148
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4062 3176 4068 3188
rect 3988 3148 4068 3176
rect 3068 3108 3096 3136
rect 3988 3117 4016 3148
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4433 3179 4491 3185
rect 4212 3148 4292 3176
rect 4212 3136 4218 3148
rect 3973 3111 4031 3117
rect 3068 3080 3832 3108
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2866 3040 2872 3052
rect 2547 3012 2872 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2866 3000 2872 3012
rect 2924 3040 2930 3052
rect 3418 3040 3424 3052
rect 2924 3012 3424 3040
rect 2924 3000 2930 3012
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 3513 3046 3571 3049
rect 3694 3046 3700 3052
rect 3513 3043 3700 3046
rect 3513 3009 3525 3043
rect 3559 3018 3700 3043
rect 3559 3009 3571 3018
rect 3513 3003 3571 3009
rect 3694 3000 3700 3018
rect 3752 3000 3758 3052
rect 3804 3046 3832 3080
rect 3973 3077 3985 3111
rect 4019 3077 4031 3111
rect 3973 3071 4031 3077
rect 3865 3049 3923 3055
rect 3865 3046 3877 3049
rect 3804 3018 3877 3046
rect 3865 3015 3877 3018
rect 3911 3015 3923 3049
rect 3865 3009 3923 3015
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 4264 3049 4292 3148
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4890 3176 4896 3188
rect 4479 3148 4896 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 5902 3176 5908 3188
rect 5675 3148 5908 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6638 3136 6644 3188
rect 6696 3136 6702 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7742 3176 7748 3188
rect 7331 3148 7748 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8110 3176 8116 3188
rect 7975 3148 8116 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8202 3136 8208 3188
rect 8260 3136 8266 3188
rect 8570 3176 8576 3188
rect 8404 3148 8576 3176
rect 5184 3108 5212 3136
rect 4356 3080 5212 3108
rect 5261 3111 5319 3117
rect 4356 3049 4384 3080
rect 5261 3077 5273 3111
rect 5307 3108 5319 3111
rect 6086 3108 6092 3120
rect 5307 3080 6092 3108
rect 5307 3077 5319 3080
rect 5261 3071 5319 3077
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 6656 3108 6684 3136
rect 7561 3111 7619 3117
rect 7561 3108 7573 3111
rect 6656 3080 7573 3108
rect 7561 3077 7573 3080
rect 7607 3077 7619 3111
rect 8220 3108 8248 3136
rect 8404 3117 8432 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9122 3176 9128 3188
rect 8803 3148 9128 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9232 3148 9628 3176
rect 7561 3071 7619 3077
rect 7760 3080 8248 3108
rect 8389 3111 8447 3117
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5166 3040 5172 3052
rect 5123 3012 5172 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 3712 2972 3740 3000
rect 4430 2972 4436 2984
rect 3712 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2972 4494 2984
rect 4908 2972 4936 3003
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5350 3000 5356 3052
rect 5408 3000 5414 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5868 3012 5917 3040
rect 5868 3000 5874 3012
rect 5905 3009 5917 3012
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6564 3012 6745 3040
rect 5721 2975 5779 2981
rect 5721 2972 5733 2975
rect 4488 2944 4936 2972
rect 5000 2944 5733 2972
rect 4488 2932 4494 2944
rect 3970 2904 3976 2916
rect 3436 2876 3976 2904
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 3326 2836 3332 2848
rect 2823 2808 3332 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 3436 2845 3464 2876
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 4525 2907 4583 2913
rect 4525 2904 4537 2907
rect 4120 2876 4537 2904
rect 4120 2864 4126 2876
rect 4525 2873 4537 2876
rect 4571 2873 4583 2907
rect 4525 2867 4583 2873
rect 4798 2864 4804 2916
rect 4856 2904 4862 2916
rect 5000 2904 5028 2944
rect 5721 2941 5733 2944
rect 5767 2941 5779 2975
rect 6012 2972 6040 3000
rect 6564 2972 6592 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 6012 2944 6592 2972
rect 6641 2975 6699 2981
rect 5721 2935 5779 2941
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7392 2972 7420 3003
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7760 3049 7788 3080
rect 8389 3077 8401 3111
rect 8435 3108 8447 3111
rect 8435 3080 9076 3108
rect 8435 3077 8447 3080
rect 8389 3071 8447 3077
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 8294 3040 8300 3052
rect 8251 3012 8300 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8478 3000 8484 3052
rect 8536 3000 8542 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8938 3040 8944 3052
rect 8619 3012 8944 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8588 2972 8616 3003
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 6687 2944 8616 2972
rect 9048 2972 9076 3080
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9232 3040 9260 3148
rect 9306 3068 9312 3120
rect 9364 3068 9370 3120
rect 9600 3108 9628 3148
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12216 3148 12265 3176
rect 12216 3136 12222 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12529 3179 12587 3185
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12710 3176 12716 3188
rect 12575 3148 12716 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 12802 3136 12808 3188
rect 12860 3136 12866 3188
rect 9600 3080 9812 3108
rect 9171 3012 9260 3040
rect 9324 3040 9352 3068
rect 9784 3052 9812 3080
rect 10410 3068 10416 3120
rect 10468 3108 10474 3120
rect 10468 3080 12388 3108
rect 10468 3068 10474 3080
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 9324 3012 9413 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 9539 3012 9573 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 9508 2972 9536 3003
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 12066 3000 12072 3052
rect 12124 3040 12130 3052
rect 12360 3049 12388 3080
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 12124 3012 12173 3040
rect 12124 3000 12130 3012
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12820 3040 12848 3136
rect 12483 3012 12848 3040
rect 12989 3043 13047 3049
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12989 3009 13001 3043
rect 13035 3040 13047 3043
rect 13446 3040 13452 3052
rect 13035 3012 13452 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 10410 2972 10416 2984
rect 9048 2944 10416 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 10928 2944 12848 2972
rect 10928 2932 10934 2944
rect 4856 2876 5028 2904
rect 4856 2864 4862 2876
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 8444 2876 9229 2904
rect 8444 2864 8450 2876
rect 9217 2873 9229 2876
rect 9263 2904 9275 2907
rect 11054 2904 11060 2916
rect 9263 2876 11060 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 12820 2913 12848 2944
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 5074 2836 5080 2848
rect 3743 2808 5080 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 5224 2808 6469 2836
rect 5224 2796 5230 2808
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 6457 2799 6515 2805
rect 1104 2746 13340 2768
rect 1104 2694 2479 2746
rect 2531 2694 2543 2746
rect 2595 2694 2607 2746
rect 2659 2694 2671 2746
rect 2723 2694 2735 2746
rect 2787 2694 5538 2746
rect 5590 2694 5602 2746
rect 5654 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 8597 2746
rect 8649 2694 8661 2746
rect 8713 2694 8725 2746
rect 8777 2694 8789 2746
rect 8841 2694 8853 2746
rect 8905 2694 11656 2746
rect 11708 2694 11720 2746
rect 11772 2694 11784 2746
rect 11836 2694 11848 2746
rect 11900 2694 11912 2746
rect 11964 2694 13340 2746
rect 1104 2672 13340 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 2866 2632 2872 2644
rect 2823 2604 2872 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4430 2632 4436 2644
rect 4387 2604 4436 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4430 2592 4436 2604
rect 4488 2632 4494 2644
rect 5166 2632 5172 2644
rect 4488 2604 5172 2632
rect 4488 2592 4494 2604
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 5994 2632 6000 2644
rect 5951 2604 6000 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6454 2592 6460 2644
rect 6512 2592 6518 2644
rect 8938 2592 8944 2644
rect 8996 2592 9002 2644
rect 10410 2592 10416 2644
rect 10468 2592 10474 2644
rect 12805 2635 12863 2641
rect 12805 2601 12817 2635
rect 12851 2632 12863 2635
rect 13078 2632 13084 2644
rect 12851 2604 13084 2632
rect 12851 2601 12863 2604
rect 12805 2595 12863 2601
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 6472 2564 6500 2592
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 6472 2536 7297 2564
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 6840 2437 6868 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11112 2468 11805 2496
rect 11112 2456 11118 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6144 2400 6745 2428
rect 6144 2388 6150 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7248 2400 7481 2428
rect 7248 2388 7254 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8812 2400 9137 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11532 2360 11560 2391
rect 11882 2360 11888 2372
rect 11532 2332 11888 2360
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12897 2363 12955 2369
rect 12897 2329 12909 2363
rect 12943 2360 12955 2363
rect 13262 2360 13268 2372
rect 12943 2332 13268 2360
rect 12943 2329 12955 2332
rect 12897 2323 12955 2329
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 1104 2202 13340 2224
rect 1104 2150 3139 2202
rect 3191 2150 3203 2202
rect 3255 2150 3267 2202
rect 3319 2150 3331 2202
rect 3383 2150 3395 2202
rect 3447 2150 6198 2202
rect 6250 2150 6262 2202
rect 6314 2150 6326 2202
rect 6378 2150 6390 2202
rect 6442 2150 6454 2202
rect 6506 2150 9257 2202
rect 9309 2150 9321 2202
rect 9373 2150 9385 2202
rect 9437 2150 9449 2202
rect 9501 2150 9513 2202
rect 9565 2150 12316 2202
rect 12368 2150 12380 2202
rect 12432 2150 12444 2202
rect 12496 2150 12508 2202
rect 12560 2150 12572 2202
rect 12624 2150 13340 2202
rect 1104 2128 13340 2150
<< via1 >>
rect 3139 14118 3191 14170
rect 3203 14118 3255 14170
rect 3267 14118 3319 14170
rect 3331 14118 3383 14170
rect 3395 14118 3447 14170
rect 6198 14118 6250 14170
rect 6262 14118 6314 14170
rect 6326 14118 6378 14170
rect 6390 14118 6442 14170
rect 6454 14118 6506 14170
rect 9257 14118 9309 14170
rect 9321 14118 9373 14170
rect 9385 14118 9437 14170
rect 9449 14118 9501 14170
rect 9513 14118 9565 14170
rect 12316 14118 12368 14170
rect 12380 14118 12432 14170
rect 12444 14118 12496 14170
rect 12508 14118 12560 14170
rect 12572 14118 12624 14170
rect 3608 14016 3660 14068
rect 10784 14016 10836 14068
rect 13268 13948 13320 14000
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 12072 13744 12124 13796
rect 2479 13574 2531 13626
rect 2543 13574 2595 13626
rect 2607 13574 2659 13626
rect 2671 13574 2723 13626
rect 2735 13574 2787 13626
rect 5538 13574 5590 13626
rect 5602 13574 5654 13626
rect 5666 13574 5718 13626
rect 5730 13574 5782 13626
rect 5794 13574 5846 13626
rect 8597 13574 8649 13626
rect 8661 13574 8713 13626
rect 8725 13574 8777 13626
rect 8789 13574 8841 13626
rect 8853 13574 8905 13626
rect 11656 13574 11708 13626
rect 11720 13574 11772 13626
rect 11784 13574 11836 13626
rect 11848 13574 11900 13626
rect 11912 13574 11964 13626
rect 6552 13336 6604 13388
rect 8024 13336 8076 13388
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7380 13268 7432 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7840 13132 7892 13184
rect 8392 13132 8444 13184
rect 11612 13268 11664 13320
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 3139 13030 3191 13082
rect 3203 13030 3255 13082
rect 3267 13030 3319 13082
rect 3331 13030 3383 13082
rect 3395 13030 3447 13082
rect 6198 13030 6250 13082
rect 6262 13030 6314 13082
rect 6326 13030 6378 13082
rect 6390 13030 6442 13082
rect 6454 13030 6506 13082
rect 9257 13030 9309 13082
rect 9321 13030 9373 13082
rect 9385 13030 9437 13082
rect 9449 13030 9501 13082
rect 9513 13030 9565 13082
rect 12316 13030 12368 13082
rect 12380 13030 12432 13082
rect 12444 13030 12496 13082
rect 12508 13030 12560 13082
rect 12572 13030 12624 13082
rect 7380 12928 7432 12980
rect 6644 12860 6696 12912
rect 5540 12724 5592 12776
rect 5908 12724 5960 12776
rect 6552 12724 6604 12776
rect 7288 12860 7340 12912
rect 8024 12860 8076 12912
rect 8484 12860 8536 12912
rect 7840 12724 7892 12776
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 9680 12792 9732 12844
rect 11428 12792 11480 12844
rect 12072 12792 12124 12844
rect 10140 12724 10192 12776
rect 9864 12656 9916 12708
rect 6000 12588 6052 12640
rect 7196 12588 7248 12640
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 10324 12588 10376 12640
rect 2479 12486 2531 12538
rect 2543 12486 2595 12538
rect 2607 12486 2659 12538
rect 2671 12486 2723 12538
rect 2735 12486 2787 12538
rect 5538 12486 5590 12538
rect 5602 12486 5654 12538
rect 5666 12486 5718 12538
rect 5730 12486 5782 12538
rect 5794 12486 5846 12538
rect 8597 12486 8649 12538
rect 8661 12486 8713 12538
rect 8725 12486 8777 12538
rect 8789 12486 8841 12538
rect 8853 12486 8905 12538
rect 11656 12486 11708 12538
rect 11720 12486 11772 12538
rect 11784 12486 11836 12538
rect 11848 12486 11900 12538
rect 11912 12486 11964 12538
rect 7472 12384 7524 12436
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 6552 12248 6604 12300
rect 6736 12180 6788 12232
rect 8484 12384 8536 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 8392 12359 8444 12368
rect 8392 12325 8401 12359
rect 8401 12325 8435 12359
rect 8435 12325 8444 12359
rect 8392 12316 8444 12325
rect 10416 12384 10468 12436
rect 11980 12384 12032 12436
rect 5908 12112 5960 12164
rect 7748 12180 7800 12232
rect 7380 12155 7432 12164
rect 7380 12121 7405 12155
rect 7405 12121 7432 12155
rect 7380 12112 7432 12121
rect 8116 12112 8168 12164
rect 8392 12112 8444 12164
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9036 12112 9088 12164
rect 9864 12180 9916 12232
rect 10140 12223 10192 12232
rect 10140 12189 10164 12223
rect 10164 12189 10192 12223
rect 10140 12180 10192 12189
rect 6000 12044 6052 12096
rect 7104 12044 7156 12096
rect 9634 12044 9686 12096
rect 9956 12044 10008 12096
rect 12072 12180 12124 12232
rect 10324 12044 10376 12096
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 3139 11942 3191 11994
rect 3203 11942 3255 11994
rect 3267 11942 3319 11994
rect 3331 11942 3383 11994
rect 3395 11942 3447 11994
rect 6198 11942 6250 11994
rect 6262 11942 6314 11994
rect 6326 11942 6378 11994
rect 6390 11942 6442 11994
rect 6454 11942 6506 11994
rect 9257 11942 9309 11994
rect 9321 11942 9373 11994
rect 9385 11942 9437 11994
rect 9449 11942 9501 11994
rect 9513 11942 9565 11994
rect 12316 11942 12368 11994
rect 12380 11942 12432 11994
rect 12444 11942 12496 11994
rect 12508 11942 12560 11994
rect 12572 11942 12624 11994
rect 5908 11704 5960 11756
rect 6552 11704 6604 11756
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 7288 11840 7340 11892
rect 9496 11840 9548 11892
rect 7104 11704 7156 11756
rect 10048 11840 10100 11892
rect 10232 11840 10284 11892
rect 5540 11636 5592 11688
rect 8392 11636 8444 11688
rect 9128 11636 9180 11688
rect 9588 11747 9640 11756
rect 9588 11713 9597 11747
rect 9597 11713 9631 11747
rect 9631 11713 9640 11747
rect 9588 11704 9640 11713
rect 9956 11704 10008 11756
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 10968 11704 11020 11756
rect 11980 11840 12032 11892
rect 4344 11500 4396 11552
rect 7196 11500 7248 11552
rect 8300 11500 8352 11552
rect 11520 11636 11572 11688
rect 10692 11500 10744 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 11428 11500 11480 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 2479 11398 2531 11450
rect 2543 11398 2595 11450
rect 2607 11398 2659 11450
rect 2671 11398 2723 11450
rect 2735 11398 2787 11450
rect 5538 11398 5590 11450
rect 5602 11398 5654 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 8597 11398 8649 11450
rect 8661 11398 8713 11450
rect 8725 11398 8777 11450
rect 8789 11398 8841 11450
rect 8853 11398 8905 11450
rect 11656 11398 11708 11450
rect 11720 11398 11772 11450
rect 11784 11398 11836 11450
rect 11848 11398 11900 11450
rect 11912 11398 11964 11450
rect 4068 11296 4120 11348
rect 6000 11296 6052 11348
rect 6644 11296 6696 11348
rect 9036 11339 9088 11348
rect 9036 11305 9045 11339
rect 9045 11305 9079 11339
rect 9079 11305 9088 11339
rect 9036 11296 9088 11305
rect 10692 11296 10744 11348
rect 11152 11339 11204 11348
rect 11152 11305 11161 11339
rect 11161 11305 11195 11339
rect 11195 11305 11204 11339
rect 11152 11296 11204 11305
rect 12256 11296 12308 11348
rect 6736 11228 6788 11280
rect 6552 11160 6604 11212
rect 10048 11228 10100 11280
rect 5080 11092 5132 11144
rect 4344 11024 4396 11076
rect 4712 11024 4764 11076
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7380 11092 7432 11144
rect 10508 11160 10560 11212
rect 8300 11067 8352 11076
rect 8300 11033 8309 11067
rect 8309 11033 8343 11067
rect 8343 11033 8352 11067
rect 8300 11024 8352 11033
rect 8392 11024 8444 11076
rect 10416 11092 10468 11144
rect 11152 11092 11204 11144
rect 11428 11228 11480 11280
rect 11336 11092 11388 11144
rect 11520 11092 11572 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 6644 10956 6696 11008
rect 9588 11024 9640 11076
rect 9956 10956 10008 11008
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 11060 10956 11112 11008
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 12072 10956 12124 11008
rect 3139 10854 3191 10906
rect 3203 10854 3255 10906
rect 3267 10854 3319 10906
rect 3331 10854 3383 10906
rect 3395 10854 3447 10906
rect 6198 10854 6250 10906
rect 6262 10854 6314 10906
rect 6326 10854 6378 10906
rect 6390 10854 6442 10906
rect 6454 10854 6506 10906
rect 9257 10854 9309 10906
rect 9321 10854 9373 10906
rect 9385 10854 9437 10906
rect 9449 10854 9501 10906
rect 9513 10854 9565 10906
rect 12316 10854 12368 10906
rect 12380 10854 12432 10906
rect 12444 10854 12496 10906
rect 12508 10854 12560 10906
rect 12572 10854 12624 10906
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 5908 10752 5960 10804
rect 4804 10616 4856 10668
rect 5448 10616 5500 10668
rect 6644 10684 6696 10736
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 7012 10616 7064 10668
rect 8392 10727 8444 10736
rect 8392 10693 8401 10727
rect 8401 10693 8435 10727
rect 8435 10693 8444 10727
rect 8392 10684 8444 10693
rect 8300 10616 8352 10668
rect 10232 10752 10284 10804
rect 10692 10795 10744 10804
rect 10692 10761 10701 10795
rect 10701 10761 10735 10795
rect 10735 10761 10744 10795
rect 10692 10752 10744 10761
rect 10968 10752 11020 10804
rect 11980 10752 12032 10804
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 12624 10684 12676 10736
rect 6552 10548 6604 10600
rect 7380 10548 7432 10600
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 6736 10480 6788 10532
rect 10600 10480 10652 10532
rect 10968 10548 11020 10600
rect 11060 10480 11112 10532
rect 11520 10616 11572 10668
rect 12072 10616 12124 10668
rect 12256 10616 12308 10668
rect 12348 10616 12400 10668
rect 11428 10548 11480 10600
rect 11612 10548 11664 10600
rect 11520 10523 11572 10532
rect 8392 10412 8444 10464
rect 9588 10412 9640 10464
rect 10968 10412 11020 10464
rect 11520 10489 11529 10523
rect 11529 10489 11563 10523
rect 11563 10489 11572 10523
rect 11520 10480 11572 10489
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 11980 10412 12032 10464
rect 2479 10310 2531 10362
rect 2543 10310 2595 10362
rect 2607 10310 2659 10362
rect 2671 10310 2723 10362
rect 2735 10310 2787 10362
rect 5538 10310 5590 10362
rect 5602 10310 5654 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 8597 10310 8649 10362
rect 8661 10310 8713 10362
rect 8725 10310 8777 10362
rect 8789 10310 8841 10362
rect 8853 10310 8905 10362
rect 11656 10310 11708 10362
rect 11720 10310 11772 10362
rect 11784 10310 11836 10362
rect 11848 10310 11900 10362
rect 11912 10310 11964 10362
rect 6552 10208 6604 10260
rect 9772 10251 9824 10260
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 10600 10208 10652 10260
rect 10968 10208 11020 10260
rect 11704 10208 11756 10260
rect 12164 10208 12216 10260
rect 10416 10140 10468 10192
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5908 10072 5960 10124
rect 3608 10004 3660 10056
rect 5908 9936 5960 9988
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 11060 10072 11112 10124
rect 11612 10072 11664 10124
rect 11980 10072 12032 10124
rect 2964 9868 3016 9920
rect 7104 9868 7156 9920
rect 9956 9868 10008 9920
rect 11244 10004 11296 10056
rect 11520 10047 11572 10056
rect 11520 10013 11530 10047
rect 11530 10013 11564 10047
rect 11564 10013 11572 10047
rect 11520 10004 11572 10013
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 11428 9868 11480 9920
rect 11888 9868 11940 9920
rect 11980 9868 12032 9920
rect 12072 9868 12124 9920
rect 12348 9868 12400 9920
rect 3139 9766 3191 9818
rect 3203 9766 3255 9818
rect 3267 9766 3319 9818
rect 3331 9766 3383 9818
rect 3395 9766 3447 9818
rect 6198 9766 6250 9818
rect 6262 9766 6314 9818
rect 6326 9766 6378 9818
rect 6390 9766 6442 9818
rect 6454 9766 6506 9818
rect 9257 9766 9309 9818
rect 9321 9766 9373 9818
rect 9385 9766 9437 9818
rect 9449 9766 9501 9818
rect 9513 9766 9565 9818
rect 12316 9766 12368 9818
rect 12380 9766 12432 9818
rect 12444 9766 12496 9818
rect 12508 9766 12560 9818
rect 12572 9766 12624 9818
rect 4804 9664 4856 9716
rect 2964 9596 3016 9648
rect 3240 9324 3292 9376
rect 3516 9324 3568 9376
rect 5908 9664 5960 9716
rect 7380 9664 7432 9716
rect 8484 9596 8536 9648
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 10508 9664 10560 9716
rect 11520 9664 11572 9716
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 8392 9460 8444 9512
rect 10876 9528 10928 9580
rect 11704 9528 11756 9580
rect 11980 9528 12032 9580
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 11336 9460 11388 9512
rect 11152 9392 11204 9444
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 7380 9367 7432 9376
rect 7380 9333 7389 9367
rect 7389 9333 7423 9367
rect 7423 9333 7432 9367
rect 7380 9324 7432 9333
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 11428 9324 11480 9376
rect 11520 9324 11572 9376
rect 11704 9324 11756 9376
rect 13084 9324 13136 9376
rect 2479 9222 2531 9274
rect 2543 9222 2595 9274
rect 2607 9222 2659 9274
rect 2671 9222 2723 9274
rect 2735 9222 2787 9274
rect 5538 9222 5590 9274
rect 5602 9222 5654 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 8597 9222 8649 9274
rect 8661 9222 8713 9274
rect 8725 9222 8777 9274
rect 8789 9222 8841 9274
rect 8853 9222 8905 9274
rect 11656 9222 11708 9274
rect 11720 9222 11772 9274
rect 11784 9222 11836 9274
rect 11848 9222 11900 9274
rect 11912 9222 11964 9274
rect 3240 9120 3292 9172
rect 5080 9120 5132 9172
rect 7380 9120 7432 9172
rect 8484 9120 8536 9172
rect 12164 9120 12216 9172
rect 4344 8984 4396 9036
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2964 8891 3016 8900
rect 2964 8857 2973 8891
rect 2973 8857 3007 8891
rect 3007 8857 3016 8891
rect 2964 8848 3016 8857
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 7104 8984 7156 9036
rect 11520 9052 11572 9104
rect 3516 8780 3568 8832
rect 4068 8823 4120 8832
rect 4068 8789 4077 8823
rect 4077 8789 4111 8823
rect 4111 8789 4120 8823
rect 4068 8780 4120 8789
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4436 8780 4488 8832
rect 5632 8848 5684 8900
rect 5724 8891 5776 8900
rect 5724 8857 5733 8891
rect 5733 8857 5767 8891
rect 5767 8857 5776 8891
rect 5724 8848 5776 8857
rect 12164 8916 12216 8968
rect 7288 8823 7340 8832
rect 7288 8789 7297 8823
rect 7297 8789 7331 8823
rect 7331 8789 7340 8823
rect 7288 8780 7340 8789
rect 8116 8780 8168 8832
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 3139 8678 3191 8730
rect 3203 8678 3255 8730
rect 3267 8678 3319 8730
rect 3331 8678 3383 8730
rect 3395 8678 3447 8730
rect 6198 8678 6250 8730
rect 6262 8678 6314 8730
rect 6326 8678 6378 8730
rect 6390 8678 6442 8730
rect 6454 8678 6506 8730
rect 9257 8678 9309 8730
rect 9321 8678 9373 8730
rect 9385 8678 9437 8730
rect 9449 8678 9501 8730
rect 9513 8678 9565 8730
rect 12316 8678 12368 8730
rect 12380 8678 12432 8730
rect 12444 8678 12496 8730
rect 12508 8678 12560 8730
rect 12572 8678 12624 8730
rect 1492 8576 1544 8628
rect 2044 8576 2096 8628
rect 2964 8576 3016 8628
rect 3608 8576 3660 8628
rect 4344 8576 4396 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 7288 8576 7340 8628
rect 10508 8576 10560 8628
rect 12164 8576 12216 8628
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3332 8440 3384 8492
rect 3884 8440 3936 8492
rect 4252 8440 4304 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 6000 8508 6052 8560
rect 3056 8372 3108 8424
rect 5632 8440 5684 8492
rect 8300 8440 8352 8492
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 4068 8304 4120 8356
rect 2228 8236 2280 8288
rect 2780 8236 2832 8288
rect 4620 8236 4672 8288
rect 7656 8279 7708 8288
rect 7656 8245 7665 8279
rect 7665 8245 7699 8279
rect 7699 8245 7708 8279
rect 7656 8236 7708 8245
rect 12440 8236 12492 8288
rect 2479 8134 2531 8186
rect 2543 8134 2595 8186
rect 2607 8134 2659 8186
rect 2671 8134 2723 8186
rect 2735 8134 2787 8186
rect 5538 8134 5590 8186
rect 5602 8134 5654 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 8597 8134 8649 8186
rect 8661 8134 8713 8186
rect 8725 8134 8777 8186
rect 8789 8134 8841 8186
rect 8853 8134 8905 8186
rect 11656 8134 11708 8186
rect 11720 8134 11772 8186
rect 11784 8134 11836 8186
rect 11848 8134 11900 8186
rect 11912 8134 11964 8186
rect 2228 8032 2280 8084
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2872 8032 2924 8084
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 4344 8032 4396 8084
rect 5080 8032 5132 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 2688 7828 2740 7880
rect 9128 7896 9180 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 7656 7828 7708 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8484 7828 8536 7880
rect 9956 7828 10008 7880
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 2320 7760 2372 7812
rect 8944 7803 8996 7812
rect 8944 7769 8953 7803
rect 8953 7769 8987 7803
rect 8987 7769 8996 7803
rect 8944 7760 8996 7769
rect 10140 7760 10192 7812
rect 12440 7760 12492 7812
rect 2228 7735 2280 7744
rect 2228 7701 2237 7735
rect 2237 7701 2271 7735
rect 2271 7701 2280 7735
rect 2228 7692 2280 7701
rect 6552 7692 6604 7744
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 9588 7692 9640 7744
rect 3139 7590 3191 7642
rect 3203 7590 3255 7642
rect 3267 7590 3319 7642
rect 3331 7590 3383 7642
rect 3395 7590 3447 7642
rect 6198 7590 6250 7642
rect 6262 7590 6314 7642
rect 6326 7590 6378 7642
rect 6390 7590 6442 7642
rect 6454 7590 6506 7642
rect 9257 7590 9309 7642
rect 9321 7590 9373 7642
rect 9385 7590 9437 7642
rect 9449 7590 9501 7642
rect 9513 7590 9565 7642
rect 12316 7590 12368 7642
rect 12380 7590 12432 7642
rect 12444 7590 12496 7642
rect 12508 7590 12560 7642
rect 12572 7590 12624 7642
rect 2412 7488 2464 7540
rect 2688 7352 2740 7404
rect 2964 7352 3016 7404
rect 3516 7352 3568 7404
rect 5908 7352 5960 7404
rect 8392 7488 8444 7540
rect 8024 7420 8076 7472
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9588 7420 9640 7472
rect 11152 7420 11204 7472
rect 9036 7352 9088 7361
rect 12072 7352 12124 7404
rect 11428 7284 11480 7336
rect 4988 7216 5040 7268
rect 4620 7148 4672 7200
rect 6000 7191 6052 7200
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 6552 7148 6604 7200
rect 6920 7148 6972 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 10140 7148 10192 7200
rect 12440 7148 12492 7200
rect 2479 7046 2531 7098
rect 2543 7046 2595 7098
rect 2607 7046 2659 7098
rect 2671 7046 2723 7098
rect 2735 7046 2787 7098
rect 5538 7046 5590 7098
rect 5602 7046 5654 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 8597 7046 8649 7098
rect 8661 7046 8713 7098
rect 8725 7046 8777 7098
rect 8789 7046 8841 7098
rect 8853 7046 8905 7098
rect 11656 7046 11708 7098
rect 11720 7046 11772 7098
rect 11784 7046 11836 7098
rect 11848 7046 11900 7098
rect 11912 7046 11964 7098
rect 2228 6944 2280 6996
rect 6000 6944 6052 6996
rect 6552 6944 6604 6996
rect 8484 6944 8536 6996
rect 9588 6944 9640 6996
rect 10968 6944 11020 6996
rect 4160 6808 4212 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3056 6740 3108 6792
rect 3516 6740 3568 6792
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 5080 6808 5132 6860
rect 5448 6808 5500 6860
rect 9956 6808 10008 6860
rect 10416 6808 10468 6860
rect 5172 6740 5224 6792
rect 6920 6740 6972 6792
rect 7288 6740 7340 6792
rect 3700 6672 3752 6724
rect 4252 6672 4304 6724
rect 4436 6672 4488 6724
rect 5356 6672 5408 6724
rect 5908 6672 5960 6724
rect 7196 6672 7248 6724
rect 8944 6740 8996 6792
rect 9036 6740 9088 6792
rect 9128 6740 9180 6792
rect 2964 6604 3016 6656
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 4712 6647 4764 6656
rect 4712 6613 4721 6647
rect 4721 6613 4755 6647
rect 4755 6613 4764 6647
rect 4712 6604 4764 6613
rect 7380 6604 7432 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 9772 6740 9824 6792
rect 9864 6740 9916 6792
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10140 6715 10192 6724
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 12440 6672 12492 6724
rect 3139 6502 3191 6554
rect 3203 6502 3255 6554
rect 3267 6502 3319 6554
rect 3331 6502 3383 6554
rect 3395 6502 3447 6554
rect 6198 6502 6250 6554
rect 6262 6502 6314 6554
rect 6326 6502 6378 6554
rect 6390 6502 6442 6554
rect 6454 6502 6506 6554
rect 9257 6502 9309 6554
rect 9321 6502 9373 6554
rect 9385 6502 9437 6554
rect 9449 6502 9501 6554
rect 9513 6502 9565 6554
rect 12316 6502 12368 6554
rect 12380 6502 12432 6554
rect 12444 6502 12496 6554
rect 12508 6502 12560 6554
rect 12572 6502 12624 6554
rect 4436 6400 4488 6452
rect 4712 6400 4764 6452
rect 4988 6400 5040 6452
rect 7196 6400 7248 6452
rect 8392 6400 8444 6452
rect 8668 6400 8720 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 9772 6400 9824 6452
rect 1400 6332 1452 6384
rect 2320 6196 2372 6248
rect 3148 6264 3200 6316
rect 3056 6196 3108 6248
rect 4252 6375 4304 6384
rect 4252 6341 4261 6375
rect 4261 6341 4295 6375
rect 4295 6341 4304 6375
rect 4252 6332 4304 6341
rect 5908 6332 5960 6384
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 4068 6196 4120 6248
rect 7288 6332 7340 6384
rect 9128 6332 9180 6384
rect 9588 6307 9640 6316
rect 4252 6196 4304 6248
rect 5264 6196 5316 6248
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 9864 6375 9916 6384
rect 9864 6341 9873 6375
rect 9873 6341 9907 6375
rect 9907 6341 9916 6375
rect 9864 6332 9916 6341
rect 10048 6400 10100 6452
rect 10600 6400 10652 6452
rect 8668 6196 8720 6248
rect 9772 6196 9824 6248
rect 10416 6332 10468 6384
rect 11980 6264 12032 6316
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 2136 6060 2188 6112
rect 2872 6060 2924 6112
rect 3976 6060 4028 6112
rect 5080 6060 5132 6112
rect 2479 5958 2531 6010
rect 2543 5958 2595 6010
rect 2607 5958 2659 6010
rect 2671 5958 2723 6010
rect 2735 5958 2787 6010
rect 5538 5958 5590 6010
rect 5602 5958 5654 6010
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 8597 5958 8649 6010
rect 8661 5958 8713 6010
rect 8725 5958 8777 6010
rect 8789 5958 8841 6010
rect 8853 5958 8905 6010
rect 11656 5958 11708 6010
rect 11720 5958 11772 6010
rect 11784 5958 11836 6010
rect 11848 5958 11900 6010
rect 11912 5958 11964 6010
rect 1400 5856 1452 5908
rect 4344 5899 4396 5908
rect 4344 5865 4353 5899
rect 4353 5865 4387 5899
rect 4387 5865 4396 5899
rect 4344 5856 4396 5865
rect 4436 5856 4488 5908
rect 4528 5856 4580 5908
rect 4896 5856 4948 5908
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 5172 5856 5224 5908
rect 6920 5856 6972 5908
rect 2136 5720 2188 5772
rect 2872 5652 2924 5704
rect 3976 5516 4028 5568
rect 8760 5788 8812 5840
rect 9036 5720 9088 5772
rect 7012 5516 7064 5568
rect 8208 5584 8260 5636
rect 3139 5414 3191 5466
rect 3203 5414 3255 5466
rect 3267 5414 3319 5466
rect 3331 5414 3383 5466
rect 3395 5414 3447 5466
rect 6198 5414 6250 5466
rect 6262 5414 6314 5466
rect 6326 5414 6378 5466
rect 6390 5414 6442 5466
rect 6454 5414 6506 5466
rect 9257 5414 9309 5466
rect 9321 5414 9373 5466
rect 9385 5414 9437 5466
rect 9449 5414 9501 5466
rect 9513 5414 9565 5466
rect 12316 5414 12368 5466
rect 12380 5414 12432 5466
rect 12444 5414 12496 5466
rect 12508 5414 12560 5466
rect 12572 5414 12624 5466
rect 3056 5312 3108 5364
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 5264 5312 5316 5364
rect 5908 5312 5960 5364
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 9128 5312 9180 5364
rect 9772 5312 9824 5364
rect 9864 5312 9916 5364
rect 2320 5244 2372 5296
rect 4068 5244 4120 5296
rect 5540 5287 5592 5296
rect 5540 5253 5549 5287
rect 5549 5253 5583 5287
rect 5583 5253 5592 5287
rect 5540 5244 5592 5253
rect 8300 5287 8352 5296
rect 8300 5253 8317 5287
rect 8317 5253 8352 5287
rect 8300 5244 8352 5253
rect 3700 5176 3752 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 6920 5176 6972 5228
rect 8300 5108 8352 5160
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 9220 5176 9272 5228
rect 10692 5287 10744 5296
rect 10692 5253 10701 5287
rect 10701 5253 10735 5287
rect 10735 5253 10744 5287
rect 10692 5244 10744 5253
rect 11060 5244 11112 5296
rect 9864 5108 9916 5160
rect 11428 5108 11480 5160
rect 2136 4972 2188 5024
rect 4344 4972 4396 5024
rect 8208 4972 8260 5024
rect 9772 4972 9824 5024
rect 11244 4972 11296 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 12164 4972 12216 5024
rect 2479 4870 2531 4922
rect 2543 4870 2595 4922
rect 2607 4870 2659 4922
rect 2671 4870 2723 4922
rect 2735 4870 2787 4922
rect 5538 4870 5590 4922
rect 5602 4870 5654 4922
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 8597 4870 8649 4922
rect 8661 4870 8713 4922
rect 8725 4870 8777 4922
rect 8789 4870 8841 4922
rect 8853 4870 8905 4922
rect 11656 4870 11708 4922
rect 11720 4870 11772 4922
rect 11784 4870 11836 4922
rect 11848 4870 11900 4922
rect 11912 4870 11964 4922
rect 9220 4768 9272 4820
rect 11428 4768 11480 4820
rect 12808 4768 12860 4820
rect 4804 4632 4856 4684
rect 11520 4632 11572 4684
rect 940 4564 992 4616
rect 2136 4428 2188 4480
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 10968 4496 11020 4548
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 12164 4496 12216 4548
rect 11060 4428 11112 4480
rect 11336 4428 11388 4480
rect 3139 4326 3191 4378
rect 3203 4326 3255 4378
rect 3267 4326 3319 4378
rect 3331 4326 3383 4378
rect 3395 4326 3447 4378
rect 6198 4326 6250 4378
rect 6262 4326 6314 4378
rect 6326 4326 6378 4378
rect 6390 4326 6442 4378
rect 6454 4326 6506 4378
rect 9257 4326 9309 4378
rect 9321 4326 9373 4378
rect 9385 4326 9437 4378
rect 9449 4326 9501 4378
rect 9513 4326 9565 4378
rect 12316 4326 12368 4378
rect 12380 4326 12432 4378
rect 12444 4326 12496 4378
rect 12508 4326 12560 4378
rect 12572 4326 12624 4378
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 4160 4267 4212 4276
rect 4160 4233 4169 4267
rect 4169 4233 4203 4267
rect 4203 4233 4212 4267
rect 4160 4224 4212 4233
rect 2044 4020 2096 4072
rect 2228 4063 2280 4072
rect 2228 4029 2237 4063
rect 2237 4029 2271 4063
rect 2271 4029 2280 4063
rect 2228 4020 2280 4029
rect 2688 4020 2740 4072
rect 4344 4088 4396 4140
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 6000 4156 6052 4208
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 7196 4224 7248 4276
rect 7288 4224 7340 4276
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 3056 3952 3108 4004
rect 3608 3952 3660 4004
rect 3976 3952 4028 4004
rect 5356 4020 5408 4072
rect 5908 4020 5960 4072
rect 6092 4020 6144 4072
rect 6460 4020 6512 4072
rect 6828 4020 6880 4072
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 8116 4088 8168 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 5264 3995 5316 4004
rect 5264 3961 5273 3995
rect 5273 3961 5307 3995
rect 5307 3961 5316 3995
rect 5264 3952 5316 3961
rect 5448 3952 5500 4004
rect 7104 3995 7156 4004
rect 7104 3961 7113 3995
rect 7113 3961 7147 3995
rect 7147 3961 7156 3995
rect 7104 3952 7156 3961
rect 7196 3952 7248 4004
rect 2872 3884 2924 3936
rect 3884 3884 3936 3936
rect 5080 3884 5132 3936
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 6644 3884 6696 3936
rect 6920 3884 6972 3936
rect 7564 3884 7616 3936
rect 10876 4224 10928 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 11336 4224 11388 4276
rect 11060 4156 11112 4208
rect 9772 4088 9824 4140
rect 9864 4088 9916 4140
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 9128 3995 9180 4004
rect 9128 3961 9137 3995
rect 9137 3961 9171 3995
rect 9171 3961 9180 3995
rect 9128 3952 9180 3961
rect 9220 3952 9272 4004
rect 8392 3884 8444 3936
rect 8484 3884 8536 3936
rect 8944 3884 8996 3936
rect 9036 3884 9088 3936
rect 10416 3952 10468 4004
rect 11244 4020 11296 4072
rect 10784 3884 10836 3936
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 2479 3782 2531 3834
rect 2543 3782 2595 3834
rect 2607 3782 2659 3834
rect 2671 3782 2723 3834
rect 2735 3782 2787 3834
rect 5538 3782 5590 3834
rect 5602 3782 5654 3834
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 8597 3782 8649 3834
rect 8661 3782 8713 3834
rect 8725 3782 8777 3834
rect 8789 3782 8841 3834
rect 8853 3782 8905 3834
rect 11656 3782 11708 3834
rect 11720 3782 11772 3834
rect 11784 3782 11836 3834
rect 11848 3782 11900 3834
rect 11912 3782 11964 3834
rect 1584 3476 1636 3528
rect 2228 3612 2280 3664
rect 2044 3544 2096 3596
rect 2872 3680 2924 3732
rect 2964 3544 3016 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3332 3612 3384 3664
rect 3608 3476 3660 3528
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 4804 3680 4856 3732
rect 5080 3680 5132 3732
rect 6828 3680 6880 3732
rect 6092 3612 6144 3664
rect 5448 3544 5500 3596
rect 6000 3544 6052 3596
rect 6920 3612 6972 3664
rect 7104 3680 7156 3732
rect 8024 3680 8076 3732
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 2044 3340 2096 3392
rect 2872 3383 2924 3392
rect 2872 3349 2881 3383
rect 2881 3349 2915 3383
rect 2915 3349 2924 3383
rect 2872 3340 2924 3349
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 5264 3476 5316 3528
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 5816 3340 5868 3392
rect 6736 3476 6788 3528
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 7288 3544 7340 3596
rect 6920 3451 6972 3460
rect 6920 3417 6929 3451
rect 6929 3417 6963 3451
rect 6963 3417 6972 3451
rect 6920 3408 6972 3417
rect 7196 3519 7248 3528
rect 7196 3485 7205 3519
rect 7205 3485 7239 3519
rect 7239 3485 7248 3519
rect 7196 3476 7248 3485
rect 7748 3544 7800 3596
rect 8484 3544 8536 3596
rect 8852 3544 8904 3596
rect 9220 3680 9272 3732
rect 10692 3680 10744 3732
rect 10876 3680 10928 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 8208 3476 8260 3528
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 8668 3476 8720 3528
rect 9036 3476 9088 3528
rect 9404 3655 9456 3664
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 9404 3612 9456 3621
rect 9588 3612 9640 3664
rect 9772 3612 9824 3664
rect 9312 3476 9364 3528
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 9680 3519 9732 3528
rect 9680 3485 9690 3519
rect 9690 3485 9724 3519
rect 9724 3485 9732 3519
rect 9680 3476 9732 3485
rect 9772 3476 9824 3528
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 8208 3340 8260 3349
rect 8300 3340 8352 3392
rect 8944 3408 8996 3460
rect 9036 3340 9088 3392
rect 9312 3340 9364 3392
rect 9404 3340 9456 3392
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 10968 3476 11020 3528
rect 11060 3340 11112 3392
rect 12716 3408 12768 3460
rect 12164 3340 12216 3392
rect 3139 3238 3191 3290
rect 3203 3238 3255 3290
rect 3267 3238 3319 3290
rect 3331 3238 3383 3290
rect 3395 3238 3447 3290
rect 6198 3238 6250 3290
rect 6262 3238 6314 3290
rect 6326 3238 6378 3290
rect 6390 3238 6442 3290
rect 6454 3238 6506 3290
rect 9257 3238 9309 3290
rect 9321 3238 9373 3290
rect 9385 3238 9437 3290
rect 9449 3238 9501 3290
rect 9513 3238 9565 3290
rect 12316 3238 12368 3290
rect 12380 3238 12432 3290
rect 12444 3238 12496 3290
rect 12508 3238 12560 3290
rect 12572 3238 12624 3290
rect 2872 3136 2924 3188
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 3332 3136 3384 3188
rect 3884 3136 3936 3188
rect 4068 3136 4120 3188
rect 4160 3136 4212 3188
rect 2872 3000 2924 3052
rect 3424 3000 3476 3052
rect 3700 3000 3752 3052
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 4896 3136 4948 3188
rect 5172 3136 5224 3188
rect 5908 3136 5960 3188
rect 6644 3136 6696 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 7748 3136 7800 3188
rect 8116 3136 8168 3188
rect 8208 3136 8260 3188
rect 6092 3111 6144 3120
rect 6092 3077 6101 3111
rect 6101 3077 6135 3111
rect 6135 3077 6144 3111
rect 6092 3068 6144 3077
rect 8576 3136 8628 3188
rect 9128 3136 9180 3188
rect 4436 2932 4488 2984
rect 5172 3000 5224 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 5816 3000 5868 3052
rect 6000 3000 6052 3052
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 3332 2796 3384 2848
rect 3976 2864 4028 2916
rect 4068 2864 4120 2916
rect 4804 2864 4856 2916
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 8300 3000 8352 3052
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 8944 3000 8996 3052
rect 9312 3068 9364 3120
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 12164 3136 12216 3188
rect 12716 3136 12768 3188
rect 12808 3136 12860 3188
rect 10416 3068 10468 3120
rect 9772 3000 9824 3052
rect 12072 3000 12124 3052
rect 13452 3000 13504 3052
rect 10416 2932 10468 2984
rect 10876 2932 10928 2984
rect 8392 2864 8444 2916
rect 11060 2864 11112 2916
rect 5080 2796 5132 2848
rect 5172 2796 5224 2848
rect 2479 2694 2531 2746
rect 2543 2694 2595 2746
rect 2607 2694 2659 2746
rect 2671 2694 2723 2746
rect 2735 2694 2787 2746
rect 5538 2694 5590 2746
rect 5602 2694 5654 2746
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 8597 2694 8649 2746
rect 8661 2694 8713 2746
rect 8725 2694 8777 2746
rect 8789 2694 8841 2746
rect 8853 2694 8905 2746
rect 11656 2694 11708 2746
rect 11720 2694 11772 2746
rect 11784 2694 11836 2746
rect 11848 2694 11900 2746
rect 11912 2694 11964 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2872 2592 2924 2644
rect 4436 2592 4488 2644
rect 5172 2592 5224 2644
rect 6000 2592 6052 2644
rect 6460 2592 6512 2644
rect 8944 2635 8996 2644
rect 8944 2601 8953 2635
rect 8953 2601 8987 2635
rect 8987 2601 8996 2635
rect 8944 2592 8996 2601
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 13084 2592 13136 2644
rect 940 2388 992 2440
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6092 2388 6144 2440
rect 11060 2456 11112 2508
rect 7196 2388 7248 2440
rect 8760 2388 8812 2440
rect 10324 2388 10376 2440
rect 11888 2320 11940 2372
rect 13268 2320 13320 2372
rect 3139 2150 3191 2202
rect 3203 2150 3255 2202
rect 3267 2150 3319 2202
rect 3331 2150 3383 2202
rect 3395 2150 3447 2202
rect 6198 2150 6250 2202
rect 6262 2150 6314 2202
rect 6326 2150 6378 2202
rect 6390 2150 6442 2202
rect 6454 2150 6506 2202
rect 9257 2150 9309 2202
rect 9321 2150 9373 2202
rect 9385 2150 9437 2202
rect 9449 2150 9501 2202
rect 9513 2150 9565 2202
rect 12316 2150 12368 2202
rect 12380 2150 12432 2202
rect 12444 2150 12496 2202
rect 12508 2150 12560 2202
rect 12572 2150 12624 2202
<< metal2 >>
rect 3606 15801 3662 16601
rect 10782 15801 10838 16601
rect 3139 14172 3447 14181
rect 3139 14170 3145 14172
rect 3201 14170 3225 14172
rect 3281 14170 3305 14172
rect 3361 14170 3385 14172
rect 3441 14170 3447 14172
rect 3201 14118 3203 14170
rect 3383 14118 3385 14170
rect 3139 14116 3145 14118
rect 3201 14116 3225 14118
rect 3281 14116 3305 14118
rect 3361 14116 3385 14118
rect 3441 14116 3447 14118
rect 3139 14107 3447 14116
rect 3620 14074 3648 15801
rect 6198 14172 6506 14181
rect 6198 14170 6204 14172
rect 6260 14170 6284 14172
rect 6340 14170 6364 14172
rect 6420 14170 6444 14172
rect 6500 14170 6506 14172
rect 6260 14118 6262 14170
rect 6442 14118 6444 14170
rect 6198 14116 6204 14118
rect 6260 14116 6284 14118
rect 6340 14116 6364 14118
rect 6420 14116 6444 14118
rect 6500 14116 6506 14118
rect 6198 14107 6506 14116
rect 9257 14172 9565 14181
rect 9257 14170 9263 14172
rect 9319 14170 9343 14172
rect 9399 14170 9423 14172
rect 9479 14170 9503 14172
rect 9559 14170 9565 14172
rect 9319 14118 9321 14170
rect 9501 14118 9503 14170
rect 9257 14116 9263 14118
rect 9319 14116 9343 14118
rect 9399 14116 9423 14118
rect 9479 14116 9503 14118
rect 9559 14116 9565 14118
rect 9257 14107 9565 14116
rect 10796 14074 10824 15801
rect 13266 14240 13322 14249
rect 12316 14172 12624 14181
rect 13266 14175 13322 14184
rect 12316 14170 12322 14172
rect 12378 14170 12402 14172
rect 12458 14170 12482 14172
rect 12538 14170 12562 14172
rect 12618 14170 12624 14172
rect 12378 14118 12380 14170
rect 12560 14118 12562 14170
rect 12316 14116 12322 14118
rect 12378 14116 12402 14118
rect 12458 14116 12482 14118
rect 12538 14116 12562 14118
rect 12618 14116 12624 14118
rect 12316 14107 12624 14116
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 13280 14006 13308 14175
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 2479 13628 2787 13637
rect 2479 13626 2485 13628
rect 2541 13626 2565 13628
rect 2621 13626 2645 13628
rect 2701 13626 2725 13628
rect 2781 13626 2787 13628
rect 2541 13574 2543 13626
rect 2723 13574 2725 13626
rect 2479 13572 2485 13574
rect 2541 13572 2565 13574
rect 2621 13572 2645 13574
rect 2701 13572 2725 13574
rect 2781 13572 2787 13574
rect 2479 13563 2787 13572
rect 3139 13084 3447 13093
rect 3139 13082 3145 13084
rect 3201 13082 3225 13084
rect 3281 13082 3305 13084
rect 3361 13082 3385 13084
rect 3441 13082 3447 13084
rect 3201 13030 3203 13082
rect 3383 13030 3385 13082
rect 3139 13028 3145 13030
rect 3201 13028 3225 13030
rect 3281 13028 3305 13030
rect 3361 13028 3385 13030
rect 3441 13028 3447 13030
rect 3139 13019 3447 13028
rect 2479 12540 2787 12549
rect 2479 12538 2485 12540
rect 2541 12538 2565 12540
rect 2621 12538 2645 12540
rect 2701 12538 2725 12540
rect 2781 12538 2787 12540
rect 2541 12486 2543 12538
rect 2723 12486 2725 12538
rect 2479 12484 2485 12486
rect 2541 12484 2565 12486
rect 2621 12484 2645 12486
rect 2701 12484 2725 12486
rect 2781 12484 2787 12486
rect 2479 12475 2787 12484
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 3139 11996 3447 12005
rect 3139 11994 3145 11996
rect 3201 11994 3225 11996
rect 3281 11994 3305 11996
rect 3361 11994 3385 11996
rect 3441 11994 3447 11996
rect 3201 11942 3203 11994
rect 3383 11942 3385 11994
rect 3139 11940 3145 11942
rect 3201 11940 3225 11942
rect 3281 11940 3305 11942
rect 3361 11940 3385 11942
rect 3441 11940 3447 11942
rect 3139 11931 3447 11940
rect 2479 11452 2787 11461
rect 2479 11450 2485 11452
rect 2541 11450 2565 11452
rect 2621 11450 2645 11452
rect 2701 11450 2725 11452
rect 2781 11450 2787 11452
rect 2541 11398 2543 11450
rect 2723 11398 2725 11450
rect 2479 11396 2485 11398
rect 2541 11396 2565 11398
rect 2621 11396 2645 11398
rect 2701 11396 2725 11398
rect 2781 11396 2787 11398
rect 2479 11387 2787 11396
rect 4080 11354 4108 12271
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3139 10908 3447 10917
rect 3139 10906 3145 10908
rect 3201 10906 3225 10908
rect 3281 10906 3305 10908
rect 3361 10906 3385 10908
rect 3441 10906 3447 10908
rect 3201 10854 3203 10906
rect 3383 10854 3385 10906
rect 3139 10852 3145 10854
rect 3201 10852 3225 10854
rect 3281 10852 3305 10854
rect 3361 10852 3385 10854
rect 3441 10852 3447 10854
rect 3139 10843 3447 10852
rect 2479 10364 2787 10373
rect 2479 10362 2485 10364
rect 2541 10362 2565 10364
rect 2621 10362 2645 10364
rect 2701 10362 2725 10364
rect 2781 10362 2787 10364
rect 2541 10310 2543 10362
rect 2723 10310 2725 10362
rect 2479 10308 2485 10310
rect 2541 10308 2565 10310
rect 2621 10308 2645 10310
rect 2701 10308 2725 10310
rect 2781 10308 2787 10310
rect 2479 10299 2787 10308
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9654 3004 9862
rect 3139 9820 3447 9829
rect 3139 9818 3145 9820
rect 3201 9818 3225 9820
rect 3281 9818 3305 9820
rect 3361 9818 3385 9820
rect 3441 9818 3447 9820
rect 3201 9766 3203 9818
rect 3383 9766 3385 9818
rect 3139 9764 3145 9766
rect 3201 9764 3225 9766
rect 3281 9764 3305 9766
rect 3361 9764 3385 9766
rect 3441 9764 3447 9766
rect 3139 9755 3447 9764
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2479 9276 2787 9285
rect 2479 9274 2485 9276
rect 2541 9274 2565 9276
rect 2621 9274 2645 9276
rect 2701 9274 2725 9276
rect 2781 9274 2787 9276
rect 2541 9222 2543 9274
rect 2723 9222 2725 9274
rect 2479 9220 2485 9222
rect 2541 9220 2565 9222
rect 2621 9220 2645 9222
rect 2701 9220 2725 9222
rect 2781 9220 2787 9222
rect 2479 9211 2787 9220
rect 3252 9178 3280 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8634 1532 8774
rect 2976 8634 3004 8842
rect 3528 8838 3556 9318
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3139 8732 3447 8741
rect 3139 8730 3145 8732
rect 3201 8730 3225 8732
rect 3281 8730 3305 8732
rect 3361 8730 3385 8732
rect 3441 8730 3447 8732
rect 3201 8678 3203 8730
rect 3383 8678 3385 8730
rect 3139 8676 3145 8678
rect 3201 8676 3225 8678
rect 3281 8676 3305 8678
rect 3361 8676 3385 8678
rect 3441 8676 3447 8678
rect 3139 8667 3447 8676
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6390 1440 6734
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1412 5914 1440 6326
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 2056 4078 2084 8570
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2516 8344 2544 8434
rect 2332 8316 2544 8344
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 8090 2268 8230
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2332 7818 2360 8316
rect 2792 8294 2820 8434
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2479 8188 2787 8197
rect 2479 8186 2485 8188
rect 2541 8186 2565 8188
rect 2621 8186 2645 8188
rect 2701 8186 2725 8188
rect 2781 8186 2787 8188
rect 2541 8134 2543 8186
rect 2723 8134 2725 8186
rect 2479 8132 2485 8134
rect 2541 8132 2565 8134
rect 2621 8132 2645 8134
rect 2701 8132 2725 8134
rect 2781 8132 2787 8134
rect 2479 8123 2787 8132
rect 2884 8090 2912 8434
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3068 8090 3096 8366
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3344 7886 3372 8434
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7002 2268 7686
rect 2424 7546 2452 7822
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2700 7410 2728 7822
rect 2976 7410 3004 7822
rect 3139 7644 3447 7653
rect 3139 7642 3145 7644
rect 3201 7642 3225 7644
rect 3281 7642 3305 7644
rect 3361 7642 3385 7644
rect 3441 7642 3447 7644
rect 3201 7590 3203 7642
rect 3383 7590 3385 7642
rect 3139 7588 3145 7590
rect 3201 7588 3225 7590
rect 3281 7588 3305 7590
rect 3361 7588 3385 7590
rect 3441 7588 3447 7590
rect 3139 7579 3447 7588
rect 3528 7410 3556 8774
rect 3620 8634 3648 9998
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 2479 7100 2787 7109
rect 2479 7098 2485 7100
rect 2541 7098 2565 7100
rect 2621 7098 2645 7100
rect 2701 7098 2725 7100
rect 2781 7098 2787 7100
rect 2541 7046 2543 7098
rect 2723 7046 2725 7098
rect 2479 7044 2485 7046
rect 2541 7044 2565 7046
rect 2621 7044 2645 7046
rect 2701 7044 2725 7046
rect 2781 7044 2787 7046
rect 2479 7035 2787 7044
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2976 6662 3004 7346
rect 3528 6798 3556 7346
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5778 2176 6054
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2332 5302 2360 6190
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2479 6012 2787 6021
rect 2479 6010 2485 6012
rect 2541 6010 2565 6012
rect 2621 6010 2645 6012
rect 2701 6010 2725 6012
rect 2781 6010 2787 6012
rect 2541 5958 2543 6010
rect 2723 5958 2725 6010
rect 2479 5956 2485 5958
rect 2541 5956 2565 5958
rect 2621 5956 2645 5958
rect 2701 5956 2725 5958
rect 2781 5956 2787 5958
rect 2479 5947 2787 5956
rect 2884 5710 2912 6054
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4486 2176 4966
rect 2479 4924 2787 4933
rect 2479 4922 2485 4924
rect 2541 4922 2565 4924
rect 2621 4922 2645 4924
rect 2701 4922 2725 4924
rect 2781 4922 2787 4924
rect 2541 4870 2543 4922
rect 2723 4870 2725 4922
rect 2479 4868 2485 4870
rect 2541 4868 2565 4870
rect 2621 4868 2645 4870
rect 2701 4868 2725 4870
rect 2781 4868 2787 4870
rect 2479 4859 2787 4868
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2228 4072 2280 4078
rect 2688 4072 2740 4078
rect 2228 4014 2280 4020
rect 2686 4040 2688 4049
rect 2740 4040 2742 4049
rect 2056 3602 2084 4014
rect 2240 3670 2268 4014
rect 2686 3975 2742 3984
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2976 3890 3004 6598
rect 3068 6440 3096 6734
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3139 6556 3447 6565
rect 3139 6554 3145 6556
rect 3201 6554 3225 6556
rect 3281 6554 3305 6556
rect 3361 6554 3385 6556
rect 3441 6554 3447 6556
rect 3201 6502 3203 6554
rect 3383 6502 3385 6554
rect 3139 6500 3145 6502
rect 3201 6500 3225 6502
rect 3281 6500 3305 6502
rect 3361 6500 3385 6502
rect 3441 6500 3447 6502
rect 3139 6491 3447 6500
rect 3068 6412 3188 6440
rect 3160 6322 3188 6412
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3712 6254 3740 6666
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3068 5370 3096 6190
rect 3139 5468 3447 5477
rect 3139 5466 3145 5468
rect 3201 5466 3225 5468
rect 3281 5466 3305 5468
rect 3361 5466 3385 5468
rect 3441 5466 3447 5468
rect 3201 5414 3203 5466
rect 3383 5414 3385 5466
rect 3139 5412 3145 5414
rect 3201 5412 3225 5414
rect 3281 5412 3305 5414
rect 3361 5412 3385 5414
rect 3441 5412 3447 5414
rect 3139 5403 3447 5412
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3712 5234 3740 6190
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3139 4380 3447 4389
rect 3139 4378 3145 4380
rect 3201 4378 3225 4380
rect 3281 4378 3305 4380
rect 3361 4378 3385 4380
rect 3441 4378 3447 4380
rect 3201 4326 3203 4378
rect 3383 4326 3385 4378
rect 3139 4324 3145 4326
rect 3201 4324 3225 4326
rect 3281 4324 3305 4326
rect 3361 4324 3385 4326
rect 3441 4324 3447 4326
rect 3139 4315 3447 4324
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 3068 3890 3096 3946
rect 2479 3836 2787 3845
rect 2479 3834 2485 3836
rect 2541 3834 2565 3836
rect 2621 3834 2645 3836
rect 2701 3834 2725 3836
rect 2781 3834 2787 3836
rect 2541 3782 2543 3834
rect 2723 3782 2725 3834
rect 2479 3780 2485 3782
rect 2541 3780 2565 3782
rect 2621 3780 2645 3782
rect 2701 3780 2725 3782
rect 2781 3780 2787 3782
rect 2479 3771 2787 3780
rect 2884 3738 2912 3878
rect 2976 3862 3096 3890
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2228 3664 2280 3670
rect 2228 3606 2280 3612
rect 2976 3602 3004 3862
rect 3344 3670 3372 4218
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 2650 1624 3470
rect 2056 3398 2084 3538
rect 3620 3534 3648 3946
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2884 3194 2912 3334
rect 3068 3194 3096 3470
rect 3139 3292 3447 3301
rect 3139 3290 3145 3292
rect 3201 3290 3225 3292
rect 3281 3290 3305 3292
rect 3361 3290 3385 3292
rect 3441 3290 3447 3292
rect 3201 3238 3203 3290
rect 3383 3238 3385 3290
rect 3139 3236 3145 3238
rect 3201 3236 3225 3238
rect 3281 3236 3305 3238
rect 3361 3236 3385 3238
rect 3441 3236 3447 3238
rect 3139 3227 3447 3236
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2479 2748 2787 2757
rect 2479 2746 2485 2748
rect 2541 2746 2565 2748
rect 2621 2746 2645 2748
rect 2701 2746 2725 2748
rect 2781 2746 2787 2748
rect 2541 2694 2543 2746
rect 2723 2694 2725 2746
rect 2479 2692 2485 2694
rect 2541 2692 2565 2694
rect 2621 2692 2645 2694
rect 2701 2692 2725 2694
rect 2781 2692 2787 2694
rect 2479 2683 2787 2692
rect 2884 2650 2912 2994
rect 3344 2854 3372 3130
rect 3620 3074 3648 3470
rect 3436 3058 3648 3074
rect 3712 3058 3740 4014
rect 3896 3942 3924 8434
rect 4080 8362 4108 8774
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 6254 4108 8298
rect 4172 6866 4200 13874
rect 5538 13628 5846 13637
rect 5538 13626 5544 13628
rect 5600 13626 5624 13628
rect 5680 13626 5704 13628
rect 5760 13626 5784 13628
rect 5840 13626 5846 13628
rect 5600 13574 5602 13626
rect 5782 13574 5784 13626
rect 5538 13572 5544 13574
rect 5600 13572 5624 13574
rect 5680 13572 5704 13574
rect 5760 13572 5784 13574
rect 5840 13572 5846 13574
rect 5538 13563 5846 13572
rect 8597 13628 8905 13637
rect 8597 13626 8603 13628
rect 8659 13626 8683 13628
rect 8739 13626 8763 13628
rect 8819 13626 8843 13628
rect 8899 13626 8905 13628
rect 8659 13574 8661 13626
rect 8841 13574 8843 13626
rect 8597 13572 8603 13574
rect 8659 13572 8683 13574
rect 8739 13572 8763 13574
rect 8819 13572 8843 13574
rect 8899 13572 8905 13574
rect 8597 13563 8905 13572
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 6198 13084 6506 13093
rect 6198 13082 6204 13084
rect 6260 13082 6284 13084
rect 6340 13082 6364 13084
rect 6420 13082 6444 13084
rect 6500 13082 6506 13084
rect 6260 13030 6262 13082
rect 6442 13030 6444 13082
rect 6198 13028 6204 13030
rect 6260 13028 6284 13030
rect 6340 13028 6364 13030
rect 6420 13028 6444 13030
rect 6500 13028 6506 13030
rect 6198 13019 6506 13028
rect 6564 12782 6592 13330
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7300 12918 7328 13262
rect 7392 12986 7420 13262
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 5552 12628 5580 12718
rect 5460 12600 5580 12628
rect 5460 12434 5488 12600
rect 5538 12540 5846 12549
rect 5538 12538 5544 12540
rect 5600 12538 5624 12540
rect 5680 12538 5704 12540
rect 5760 12538 5784 12540
rect 5840 12538 5846 12540
rect 5600 12486 5602 12538
rect 5782 12486 5784 12538
rect 5538 12484 5544 12486
rect 5600 12484 5624 12486
rect 5680 12484 5704 12486
rect 5760 12484 5784 12486
rect 5840 12484 5846 12486
rect 5538 12475 5846 12484
rect 5460 12406 5580 12434
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11082 4384 11494
rect 5092 11150 5120 12242
rect 5552 11694 5580 12406
rect 5920 12170 5948 12718
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 6012 12102 6040 12582
rect 6564 12306 6592 12718
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6198 11996 6506 12005
rect 6198 11994 6204 11996
rect 6260 11994 6284 11996
rect 6340 11994 6364 11996
rect 6420 11994 6444 11996
rect 6500 11994 6506 11996
rect 6260 11942 6262 11994
rect 6442 11942 6444 11994
rect 6198 11940 6204 11942
rect 6260 11940 6284 11942
rect 6340 11940 6364 11942
rect 6420 11940 6444 11942
rect 6500 11940 6506 11942
rect 6198 11931 6506 11940
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 5540 11688 5592 11694
rect 5460 11636 5540 11642
rect 5460 11630 5592 11636
rect 5460 11614 5580 11630
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4724 10810 4752 11018
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 9722 4844 10610
rect 5092 10130 5120 11086
rect 5460 10674 5488 11614
rect 5538 11452 5846 11461
rect 5538 11450 5544 11452
rect 5600 11450 5624 11452
rect 5680 11450 5704 11452
rect 5760 11450 5784 11452
rect 5840 11450 5846 11452
rect 5600 11398 5602 11450
rect 5782 11398 5784 11450
rect 5538 11396 5544 11398
rect 5600 11396 5624 11398
rect 5680 11396 5704 11398
rect 5760 11396 5784 11398
rect 5840 11396 5846 11398
rect 5538 11387 5846 11396
rect 5920 10810 5948 11698
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5538 10364 5846 10373
rect 5538 10362 5544 10364
rect 5600 10362 5624 10364
rect 5680 10362 5704 10364
rect 5760 10362 5784 10364
rect 5840 10362 5846 10364
rect 5600 10310 5602 10362
rect 5782 10310 5784 10362
rect 5538 10308 5544 10310
rect 5600 10308 5624 10310
rect 5680 10308 5704 10310
rect 5760 10308 5784 10310
rect 5840 10308 5846 10310
rect 5538 10299 5846 10308
rect 5920 10130 5948 10406
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 9042 4384 9318
rect 4344 9036 4396 9042
rect 4264 8996 4344 9024
rect 4264 8498 4292 8996
rect 4344 8978 4396 8984
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4356 8634 4384 8774
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4448 8514 4476 8774
rect 4356 8498 4476 8514
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4344 8492 4476 8498
rect 4396 8486 4476 8492
rect 4344 8434 4396 8440
rect 4356 8090 4384 8434
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4632 7206 4660 8230
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4264 6390 4292 6666
rect 4448 6458 4476 6666
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4264 6254 4292 6326
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5574 4016 6054
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 5234 4016 5510
rect 4080 5302 4108 6190
rect 4448 5914 4476 6394
rect 4540 5914 4568 6598
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4356 5794 4384 5850
rect 4632 5794 4660 7142
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 6458 4752 6598
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4356 5766 4660 5794
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 4010 4016 5170
rect 4356 5030 4384 5766
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4816 4690 4844 9658
rect 5092 9178 5120 10066
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5920 9722 5948 9930
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5538 9276 5846 9285
rect 5538 9274 5544 9276
rect 5600 9274 5624 9276
rect 5680 9274 5704 9276
rect 5760 9274 5784 9276
rect 5840 9274 5846 9276
rect 5600 9222 5602 9274
rect 5782 9222 5784 9274
rect 5538 9220 5544 9222
rect 5600 9220 5624 9222
rect 5680 9220 5704 9222
rect 5760 9220 5784 9222
rect 5840 9220 5846 9222
rect 5538 9211 5846 9220
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5092 8090 5120 9114
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 5914 4936 6734
rect 5000 6458 5028 7210
rect 5460 6866 5488 8910
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5644 8498 5672 8842
rect 5736 8634 5764 8842
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 6012 8566 6040 11290
rect 6564 11218 6592 11698
rect 6656 11354 6684 12854
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6748 11286 6776 12174
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11762 7144 12038
rect 7208 11898 7236 12582
rect 7300 11898 7328 12854
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12170 7420 12582
rect 7484 12442 7512 13126
rect 7852 12782 7880 13126
rect 8036 12918 8064 13330
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7472 12436 7524 12442
rect 8036 12434 8064 12854
rect 7472 12378 7524 12384
rect 7760 12406 8064 12434
rect 7760 12238 7788 12406
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11642 7144 11698
rect 7116 11614 7328 11642
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6198 10908 6506 10917
rect 6198 10906 6204 10908
rect 6260 10906 6284 10908
rect 6340 10906 6364 10908
rect 6420 10906 6444 10908
rect 6500 10906 6506 10908
rect 6260 10854 6262 10906
rect 6442 10854 6444 10906
rect 6198 10852 6204 10854
rect 6260 10852 6284 10854
rect 6340 10852 6364 10854
rect 6420 10852 6444 10854
rect 6500 10852 6506 10854
rect 6198 10843 6506 10852
rect 6564 10606 6592 11154
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10742 6684 10950
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 10266 6592 10542
rect 6748 10538 6776 11222
rect 7208 11150 7236 11494
rect 7300 11150 7328 11614
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7024 10674 7052 11086
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 7024 10010 7052 10610
rect 7392 10606 7420 11086
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 10062 7420 10542
rect 7380 10056 7432 10062
rect 7024 9982 7144 10010
rect 7380 9998 7432 10004
rect 7116 9926 7144 9982
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6198 9820 6506 9829
rect 6198 9818 6204 9820
rect 6260 9818 6284 9820
rect 6340 9818 6364 9820
rect 6420 9818 6444 9820
rect 6500 9818 6506 9820
rect 6260 9766 6262 9818
rect 6442 9766 6444 9818
rect 6198 9764 6204 9766
rect 6260 9764 6284 9766
rect 6340 9764 6364 9766
rect 6420 9764 6444 9766
rect 6500 9764 6506 9766
rect 6198 9755 6506 9764
rect 7116 9042 7144 9862
rect 7392 9722 7420 9998
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7760 9586 7788 12174
rect 8128 12170 8156 13262
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12374 8432 13126
rect 9257 13084 9565 13093
rect 9257 13082 9263 13084
rect 9319 13082 9343 13084
rect 9399 13082 9423 13084
rect 9479 13082 9503 13084
rect 9559 13082 9565 13084
rect 9319 13030 9321 13082
rect 9501 13030 9503 13082
rect 9257 13028 9263 13030
rect 9319 13028 9343 13030
rect 9399 13028 9423 13030
rect 9479 13028 9503 13030
rect 9559 13028 9565 13030
rect 9257 13019 9565 13028
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8496 12442 8524 12854
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 8597 12540 8905 12549
rect 8597 12538 8603 12540
rect 8659 12538 8683 12540
rect 8739 12538 8763 12540
rect 8819 12538 8843 12540
rect 8899 12538 8905 12540
rect 8659 12486 8661 12538
rect 8841 12486 8843 12538
rect 8597 12484 8603 12486
rect 8659 12484 8683 12486
rect 8739 12484 8763 12486
rect 8819 12484 8843 12486
rect 8899 12484 8905 12486
rect 8597 12475 8905 12484
rect 9692 12442 9720 12786
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 9876 12238 9904 12650
rect 10152 12238 10180 12718
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 9128 12232 9180 12238
rect 8390 12200 8446 12209
rect 8116 12164 8168 12170
rect 9864 12232 9916 12238
rect 9128 12174 9180 12180
rect 9784 12192 9864 12220
rect 8390 12135 8392 12144
rect 8116 12106 8168 12112
rect 8444 12135 8446 12144
rect 9036 12164 9088 12170
rect 8392 12106 8444 12112
rect 9036 12106 9088 12112
rect 8404 11694 8432 12106
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 11082 8340 11494
rect 8597 11452 8905 11461
rect 8597 11450 8603 11452
rect 8659 11450 8683 11452
rect 8739 11450 8763 11452
rect 8819 11450 8843 11452
rect 8899 11450 8905 11452
rect 8659 11398 8661 11450
rect 8841 11398 8843 11450
rect 8597 11396 8603 11398
rect 8659 11396 8683 11398
rect 8739 11396 8763 11398
rect 8819 11396 8843 11398
rect 8899 11396 8905 11398
rect 8597 11387 8905 11396
rect 9048 11354 9076 12106
rect 9140 11694 9168 12174
rect 9634 12096 9686 12102
rect 9686 12064 9734 12073
rect 9634 12038 9678 12044
rect 9646 12022 9678 12038
rect 9257 11996 9565 12005
rect 9678 11999 9734 12008
rect 9257 11994 9263 11996
rect 9319 11994 9343 11996
rect 9399 11994 9423 11996
rect 9479 11994 9503 11996
rect 9559 11994 9565 11996
rect 9319 11942 9321 11994
rect 9501 11942 9503 11994
rect 9257 11940 9263 11942
rect 9319 11940 9343 11942
rect 9399 11940 9423 11942
rect 9479 11940 9503 11942
rect 9559 11940 9565 11942
rect 9257 11931 9565 11940
rect 9784 11914 9812 12192
rect 9864 12174 9916 12180
rect 10140 12232 10192 12238
rect 10192 12192 10272 12220
rect 10140 12174 10192 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 10138 12064 10194 12073
rect 9496 11892 9548 11898
rect 9600 11886 9812 11914
rect 9600 11880 9628 11886
rect 9548 11852 9628 11880
rect 9496 11834 9548 11840
rect 9968 11762 9996 12038
rect 10138 11999 10194 12008
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9600 11082 9628 11698
rect 10060 11286 10088 11834
rect 10152 11762 10180 11999
rect 10244 11898 10272 12192
rect 10336 12102 10364 12582
rect 10416 12436 10468 12442
rect 10980 12434 11008 13874
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 11656 13628 11964 13637
rect 11656 13626 11662 13628
rect 11718 13626 11742 13628
rect 11798 13626 11822 13628
rect 11878 13626 11902 13628
rect 11958 13626 11964 13628
rect 11718 13574 11720 13626
rect 11900 13574 11902 13626
rect 11656 13572 11662 13574
rect 11718 13572 11742 13574
rect 11798 13572 11822 13574
rect 11878 13572 11902 13574
rect 11958 13572 11964 13574
rect 11656 13563 11964 13572
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12986 11652 13262
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11440 12434 11468 12786
rect 11656 12540 11964 12549
rect 11656 12538 11662 12540
rect 11718 12538 11742 12540
rect 11798 12538 11822 12540
rect 11878 12538 11902 12540
rect 11958 12538 11964 12540
rect 11718 12486 11720 12538
rect 11900 12486 11902 12538
rect 11656 12484 11662 12486
rect 11718 12484 11742 12486
rect 11798 12484 11822 12486
rect 11878 12484 11902 12486
rect 11958 12484 11964 12486
rect 11656 12475 11964 12484
rect 11992 12442 12020 13126
rect 12084 12850 12112 13738
rect 12316 13084 12624 13093
rect 12316 13082 12322 13084
rect 12378 13082 12402 13084
rect 12458 13082 12482 13084
rect 12538 13082 12562 13084
rect 12618 13082 12624 13084
rect 12378 13030 12380 13082
rect 12560 13030 12562 13082
rect 12316 13028 12322 13030
rect 12378 13028 12402 13030
rect 12458 13028 12482 13030
rect 12538 13028 12562 13030
rect 12618 13028 12624 13030
rect 12316 13019 12624 13028
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 10416 12378 10468 12384
rect 10888 12406 11008 12434
rect 11072 12406 11468 12434
rect 11980 12436 12032 12442
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10232 11892 10284 11898
rect 10428 11880 10456 12378
rect 10232 11834 10284 11840
rect 10336 11852 10456 11880
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10336 11336 10364 11852
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10244 11308 10364 11336
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 8312 10674 8340 11018
rect 8404 10742 8432 11018
rect 9257 10908 9565 10917
rect 9257 10906 9263 10908
rect 9319 10906 9343 10908
rect 9399 10906 9423 10908
rect 9479 10906 9503 10908
rect 9559 10906 9565 10908
rect 9319 10854 9321 10906
rect 9501 10854 9503 10906
rect 9257 10852 9263 10854
rect 9319 10852 9343 10854
rect 9399 10852 9423 10854
rect 9479 10852 9503 10854
rect 9559 10852 9565 10854
rect 9257 10843 9565 10852
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9178 7420 9318
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6198 8732 6506 8741
rect 6198 8730 6204 8732
rect 6260 8730 6284 8732
rect 6340 8730 6364 8732
rect 6420 8730 6444 8732
rect 6500 8730 6506 8732
rect 6260 8678 6262 8730
rect 6442 8678 6444 8730
rect 6198 8676 6204 8678
rect 6260 8676 6284 8678
rect 6340 8676 6364 8678
rect 6420 8676 6444 8678
rect 6500 8676 6506 8678
rect 6198 8667 6506 8676
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5538 8188 5846 8197
rect 5538 8186 5544 8188
rect 5600 8186 5624 8188
rect 5680 8186 5704 8188
rect 5760 8186 5784 8188
rect 5840 8186 5846 8188
rect 5600 8134 5602 8186
rect 5782 8134 5784 8186
rect 5538 8132 5544 8134
rect 5600 8132 5624 8134
rect 5680 8132 5704 8134
rect 5760 8132 5784 8134
rect 5840 8132 5846 8134
rect 5538 8123 5846 8132
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6198 7644 6506 7653
rect 6198 7642 6204 7644
rect 6260 7642 6284 7644
rect 6340 7642 6364 7644
rect 6420 7642 6444 7644
rect 6500 7642 6506 7644
rect 6260 7590 6262 7642
rect 6442 7590 6444 7642
rect 6198 7588 6204 7590
rect 6260 7588 6284 7590
rect 6340 7588 6364 7590
rect 6420 7588 6444 7590
rect 6500 7588 6506 7590
rect 6198 7579 6506 7588
rect 6564 7410 6592 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 5538 7100 5846 7109
rect 5538 7098 5544 7100
rect 5600 7098 5624 7100
rect 5680 7098 5704 7100
rect 5760 7098 5784 7100
rect 5840 7098 5846 7100
rect 5600 7046 5602 7098
rect 5782 7046 5784 7098
rect 5538 7044 5544 7046
rect 5600 7044 5624 7046
rect 5680 7044 5704 7046
rect 5760 7044 5784 7046
rect 5840 7044 5846 7046
rect 5538 7035 5846 7044
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5370 5028 6394
rect 5092 6118 5120 6802
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5914 5120 6054
rect 5184 5914 5212 6734
rect 5920 6730 5948 7346
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6012 7002 6040 7142
rect 6564 7002 6592 7142
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6932 6798 6960 7142
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5276 5370 5304 6190
rect 5368 5522 5396 6666
rect 6198 6556 6506 6565
rect 6198 6554 6204 6556
rect 6260 6554 6284 6556
rect 6340 6554 6364 6556
rect 6420 6554 6444 6556
rect 6500 6554 6506 6556
rect 6260 6502 6262 6554
rect 6442 6502 6444 6554
rect 6198 6500 6204 6502
rect 6260 6500 6284 6502
rect 6340 6500 6364 6502
rect 6420 6500 6444 6502
rect 6500 6500 6506 6502
rect 6198 6491 6506 6500
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5538 6012 5846 6021
rect 5538 6010 5544 6012
rect 5600 6010 5624 6012
rect 5680 6010 5704 6012
rect 5760 6010 5784 6012
rect 5840 6010 5846 6012
rect 5600 5958 5602 6010
rect 5782 5958 5784 6010
rect 5538 5956 5544 5958
rect 5600 5956 5624 5958
rect 5680 5956 5704 5958
rect 5760 5956 5784 5958
rect 5840 5956 5846 5958
rect 5538 5947 5846 5956
rect 5368 5494 5580 5522
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3194 3924 3878
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3424 3052 3648 3058
rect 3476 3046 3648 3052
rect 3700 3052 3752 3058
rect 3424 2994 3476 3000
rect 3700 2994 3752 3000
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3896 2802 3924 3130
rect 3988 2922 4016 3946
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3194 4108 3538
rect 4172 3194 4200 4218
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4356 3534 4384 4082
rect 4816 3738 4844 4082
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4080 2922 4108 2994
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4080 2802 4108 2858
rect 3896 2774 4108 2802
rect 4448 2650 4476 2926
rect 4816 2922 4844 3470
rect 4908 3194 4936 4082
rect 5276 4010 5304 5306
rect 5552 5302 5580 5494
rect 5920 5370 5948 6326
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6198 5468 6506 5477
rect 6198 5466 6204 5468
rect 6260 5466 6284 5468
rect 6340 5466 6364 5468
rect 6420 5466 6444 5468
rect 6500 5466 6506 5468
rect 6260 5414 6262 5466
rect 6442 5414 6444 5466
rect 6198 5412 6204 5414
rect 6260 5412 6284 5414
rect 6340 5412 6364 5414
rect 6420 5412 6444 5414
rect 6500 5412 6506 5414
rect 6198 5403 6506 5412
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 6932 5234 6960 5850
rect 7024 5574 7052 7822
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 5538 4924 5846 4933
rect 5538 4922 5544 4924
rect 5600 4922 5624 4924
rect 5680 4922 5704 4924
rect 5760 4922 5784 4924
rect 5840 4922 5846 4924
rect 5600 4870 5602 4922
rect 5782 4870 5784 4922
rect 5538 4868 5544 4870
rect 5600 4868 5624 4870
rect 5680 4868 5704 4870
rect 5760 4868 5784 4870
rect 5840 4868 5846 4870
rect 5538 4859 5846 4868
rect 6198 4380 6506 4389
rect 6198 4378 6204 4380
rect 6260 4378 6284 4380
rect 6340 4378 6364 4380
rect 6420 4378 6444 4380
rect 6500 4378 6506 4380
rect 6260 4326 6262 4378
rect 6442 4326 6444 4378
rect 6198 4324 6204 4326
rect 6260 4324 6284 4326
rect 6340 4324 6364 4326
rect 6420 4324 6444 4326
rect 6500 4324 6506 4326
rect 6198 4315 6506 4324
rect 7116 4264 7144 8978
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7300 8634 7328 8774
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7886 7696 8230
rect 8128 7886 8156 8774
rect 8312 8498 8340 10610
rect 9600 10470 9628 11018
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 8404 9518 8432 10406
rect 8597 10364 8905 10373
rect 8597 10362 8603 10364
rect 8659 10362 8683 10364
rect 8739 10362 8763 10364
rect 8819 10362 8843 10364
rect 8899 10362 8905 10364
rect 8659 10310 8661 10362
rect 8841 10310 8843 10362
rect 8597 10308 8603 10310
rect 8659 10308 8683 10310
rect 8739 10308 8763 10310
rect 8819 10308 8843 10310
rect 8899 10308 8905 10310
rect 8597 10299 8905 10308
rect 9784 10266 9812 10610
rect 9968 10266 9996 10950
rect 10244 10810 10272 11308
rect 10428 11150 10456 11698
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 11354 10732 11494
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9257 9820 9565 9829
rect 9257 9818 9263 9820
rect 9319 9818 9343 9820
rect 9399 9818 9423 9820
rect 9479 9818 9503 9820
rect 9559 9818 9565 9820
rect 9319 9766 9321 9818
rect 9501 9766 9503 9818
rect 9257 9764 9263 9766
rect 9319 9764 9343 9766
rect 9399 9764 9423 9766
rect 9479 9764 9503 9766
rect 9559 9764 9565 9766
rect 9257 9755 9565 9764
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8496 9178 8524 9590
rect 9784 9586 9812 10202
rect 10428 10198 10456 10610
rect 10520 10266 10548 11154
rect 10704 10810 10732 11290
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 10266 10640 10474
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9968 9518 9996 9862
rect 10520 9722 10548 10202
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10888 9586 10916 12406
rect 11072 12209 11100 12406
rect 11980 12378 12032 12384
rect 11058 12200 11114 12209
rect 11058 12135 11114 12144
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 10810 11008 11698
rect 11532 11694 11560 12038
rect 11992 11898 12020 12378
rect 12084 12238 12112 12786
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11164 11354 11192 11494
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10980 10606 11008 10746
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11072 10538 11100 10950
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10266 11008 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 11072 9382 11100 10066
rect 11164 9450 11192 11086
rect 11256 10062 11284 11494
rect 11440 11286 11468 11494
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11532 11150 11560 11630
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11656 11452 11964 11461
rect 11656 11450 11662 11452
rect 11718 11450 11742 11452
rect 11798 11450 11822 11452
rect 11878 11450 11902 11452
rect 11958 11450 11964 11452
rect 11718 11398 11720 11450
rect 11900 11398 11902 11450
rect 11656 11396 11662 11398
rect 11718 11396 11742 11398
rect 11798 11396 11822 11398
rect 11878 11396 11902 11398
rect 11958 11396 11964 11398
rect 11656 11387 11964 11396
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11348 9518 11376 11086
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10674 11560 10950
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11624 10606 11652 11086
rect 11992 10810 12020 11494
rect 12084 11150 12112 12174
rect 12316 11996 12624 12005
rect 12316 11994 12322 11996
rect 12378 11994 12402 11996
rect 12458 11994 12482 11996
rect 12538 11994 12562 11996
rect 12618 11994 12624 11996
rect 12378 11942 12380 11994
rect 12560 11942 12562 11994
rect 12316 11940 12322 11942
rect 12378 11940 12402 11942
rect 12458 11940 12482 11942
rect 12538 11940 12562 11942
rect 12618 11940 12624 11942
rect 12316 11931 12624 11940
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12268 11354 12296 11494
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11992 10554 12020 10746
rect 12084 10674 12112 10950
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11440 9926 11468 10542
rect 11520 10532 11572 10538
rect 11992 10526 12112 10554
rect 11520 10474 11572 10480
rect 11532 10146 11560 10474
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11656 10364 11964 10373
rect 11656 10362 11662 10364
rect 11718 10362 11742 10364
rect 11798 10362 11822 10364
rect 11878 10362 11902 10364
rect 11958 10362 11964 10364
rect 11718 10310 11720 10362
rect 11900 10310 11902 10362
rect 11656 10308 11662 10310
rect 11718 10308 11742 10310
rect 11798 10308 11822 10310
rect 11878 10308 11902 10310
rect 11958 10308 11964 10310
rect 11656 10299 11964 10308
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11532 10130 11652 10146
rect 11532 10124 11664 10130
rect 11532 10118 11612 10124
rect 11612 10066 11664 10072
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11716 9586 11744 10202
rect 11992 10130 12020 10406
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12084 10010 12112 10526
rect 12176 10266 12204 11086
rect 12316 10908 12624 10917
rect 12316 10906 12322 10908
rect 12378 10906 12402 10908
rect 12458 10906 12482 10908
rect 12538 10906 12562 10908
rect 12618 10906 12624 10908
rect 12378 10854 12380 10906
rect 12560 10854 12562 10906
rect 12316 10852 12322 10854
rect 12378 10852 12402 10854
rect 12458 10852 12482 10854
rect 12538 10852 12562 10854
rect 12618 10852 12624 10854
rect 12316 10843 12624 10852
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12268 10146 12296 10610
rect 11900 9982 12112 10010
rect 12176 10118 12296 10146
rect 11900 9926 11928 9982
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11992 9586 12020 9862
rect 12084 9586 12112 9862
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11440 9438 11744 9466
rect 11440 9382 11468 9438
rect 11716 9382 11744 9438
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 8597 9276 8905 9285
rect 8597 9274 8603 9276
rect 8659 9274 8683 9276
rect 8739 9274 8763 9276
rect 8819 9274 8843 9276
rect 8899 9274 8905 9276
rect 8659 9222 8661 9274
rect 8841 9222 8843 9274
rect 8597 9220 8603 9222
rect 8659 9220 8683 9222
rect 8739 9220 8763 9222
rect 8819 9220 8843 9222
rect 8899 9220 8905 9222
rect 8597 9211 8905 9220
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 9257 8732 9565 8741
rect 9257 8730 9263 8732
rect 9319 8730 9343 8732
rect 9399 8730 9423 8732
rect 9479 8730 9503 8732
rect 9559 8730 9565 8732
rect 9319 8678 9321 8730
rect 9501 8678 9503 8730
rect 9257 8676 9263 8678
rect 9319 8676 9343 8678
rect 9399 8676 9423 8678
rect 9479 8676 9503 8678
rect 9559 8676 9565 8678
rect 9257 8667 9565 8676
rect 10520 8634 10548 9318
rect 11532 9110 11560 9318
rect 11656 9276 11964 9285
rect 11656 9274 11662 9276
rect 11718 9274 11742 9276
rect 11798 9274 11822 9276
rect 11878 9274 11902 9276
rect 11958 9274 11964 9276
rect 11718 9222 11720 9274
rect 11900 9222 11902 9274
rect 11656 9220 11662 9222
rect 11718 9220 11742 9222
rect 11798 9220 11822 9222
rect 11878 9220 11902 9222
rect 11958 9220 11964 9222
rect 11656 9211 11964 9220
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7300 6798 7328 7142
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 6458 7236 6666
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7300 6390 7328 6734
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7300 4282 7328 6326
rect 7196 4276 7248 4282
rect 7116 4236 7196 4264
rect 7196 4218 7248 4224
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 6000 4208 6052 4214
rect 7392 4162 7420 6598
rect 8128 5658 8156 7822
rect 8128 5642 8248 5658
rect 8128 5636 8260 5642
rect 8128 5630 8208 5636
rect 8208 5578 8260 5584
rect 8312 5302 8340 8434
rect 8597 8188 8905 8197
rect 8597 8186 8603 8188
rect 8659 8186 8683 8188
rect 8739 8186 8763 8188
rect 8819 8186 8843 8188
rect 8899 8186 8905 8188
rect 8659 8134 8661 8186
rect 8841 8134 8843 8186
rect 8597 8132 8603 8134
rect 8659 8132 8683 8134
rect 8739 8132 8763 8134
rect 8819 8132 8843 8134
rect 8899 8132 8905 8134
rect 8597 8123 8905 8132
rect 11440 7954 11468 8774
rect 11656 8188 11964 8197
rect 11656 8186 11662 8188
rect 11718 8186 11742 8188
rect 11798 8186 11822 8188
rect 11878 8186 11902 8188
rect 11958 8186 11964 8188
rect 11718 8134 11720 8186
rect 11900 8134 11902 8186
rect 11656 8132 11662 8134
rect 11718 8132 11742 8134
rect 11798 8132 11822 8134
rect 11878 8132 11902 8134
rect 11958 8132 11964 8134
rect 11656 8123 11964 8132
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7546 8432 7686
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7002 8524 7822
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8597 7100 8905 7109
rect 8597 7098 8603 7100
rect 8659 7098 8683 7100
rect 8739 7098 8763 7100
rect 8819 7098 8843 7100
rect 8899 7098 8905 7100
rect 8659 7046 8661 7098
rect 8841 7046 8843 7098
rect 8597 7044 8603 7046
rect 8659 7044 8683 7046
rect 8739 7044 8763 7046
rect 8819 7044 8843 7046
rect 8899 7044 8905 7046
rect 8597 7035 8905 7044
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8956 6798 8984 7754
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 6798 9076 7346
rect 9140 6798 9168 7890
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9257 7644 9565 7653
rect 9257 7642 9263 7644
rect 9319 7642 9343 7644
rect 9399 7642 9423 7644
rect 9479 7642 9503 7644
rect 9559 7642 9565 7644
rect 9319 7590 9321 7642
rect 9501 7590 9503 7642
rect 9257 7588 9263 7590
rect 9319 7588 9343 7590
rect 9399 7588 9423 7590
rect 9479 7588 9503 7590
rect 9559 7588 9565 7590
rect 9257 7579 9565 7588
rect 9600 7478 9628 7686
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6458 8432 6598
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8680 6254 8708 6394
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8597 6012 8905 6021
rect 8597 6010 8603 6012
rect 8659 6010 8683 6012
rect 8739 6010 8763 6012
rect 8819 6010 8843 6012
rect 8899 6010 8905 6012
rect 8659 5958 8661 6010
rect 8841 5958 8843 6010
rect 8597 5956 8603 5958
rect 8659 5956 8683 5958
rect 8739 5956 8763 5958
rect 8819 5956 8843 5958
rect 8899 5956 8905 5958
rect 8597 5947 8905 5956
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8772 5370 8800 5782
rect 9048 5778 9076 6734
rect 9257 6556 9565 6565
rect 9257 6554 9263 6556
rect 9319 6554 9343 6556
rect 9399 6554 9423 6556
rect 9479 6554 9503 6556
rect 9559 6554 9565 6556
rect 9319 6502 9321 6554
rect 9501 6502 9503 6554
rect 9257 6500 9263 6502
rect 9319 6500 9343 6502
rect 9399 6500 9423 6502
rect 9479 6500 9503 6502
rect 9559 6500 9565 6502
rect 9257 6491 9565 6500
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9140 5370 9168 6326
rect 9600 6322 9628 6938
rect 9968 6866 9996 7822
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7206 10180 7754
rect 11164 7478 11192 7822
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9772 6792 9824 6798
rect 9692 6740 9772 6746
rect 9692 6734 9824 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9692 6718 9812 6734
rect 9692 6458 9720 6718
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6458 9812 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9876 6390 9904 6734
rect 10152 6730 10180 7142
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10140 6724 10192 6730
rect 10060 6684 10140 6712
rect 10060 6458 10088 6684
rect 10140 6666 10192 6672
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10428 6390 10456 6802
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9257 5468 9565 5477
rect 9257 5466 9263 5468
rect 9319 5466 9343 5468
rect 9399 5466 9423 5468
rect 9479 5466 9503 5468
rect 9559 5466 9565 5468
rect 9319 5414 9321 5466
rect 9501 5414 9503 5466
rect 9257 5412 9263 5414
rect 9319 5412 9343 5414
rect 9399 5412 9423 5414
rect 9479 5412 9503 5414
rect 9559 5412 9565 5414
rect 9257 5403 9565 5412
rect 9784 5370 9812 6190
rect 9876 5370 9904 6326
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10980 5250 11008 6938
rect 11164 6798 11192 7414
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 5296 11112 5302
rect 10980 5244 11060 5250
rect 10980 5238 11112 5244
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 6000 4150 6052 4156
rect 5356 4072 5408 4078
rect 5908 4072 5960 4078
rect 5356 4014 5408 4020
rect 5446 4040 5502 4049
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5092 3738 5120 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 5092 2854 5120 3470
rect 5184 3194 5212 3878
rect 5276 3534 5304 3946
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5172 3052 5224 3058
rect 5276 3040 5304 3470
rect 5368 3058 5396 4014
rect 5908 4014 5960 4020
rect 5446 3975 5448 3984
rect 5500 3975 5502 3984
rect 5448 3946 5500 3952
rect 5538 3836 5846 3845
rect 5538 3834 5544 3836
rect 5600 3834 5624 3836
rect 5680 3834 5704 3836
rect 5760 3834 5784 3836
rect 5840 3834 5846 3836
rect 5600 3782 5602 3834
rect 5782 3782 5784 3834
rect 5538 3780 5544 3782
rect 5600 3780 5624 3782
rect 5680 3780 5704 3782
rect 5760 3780 5784 3782
rect 5840 3780 5846 3782
rect 5538 3771 5846 3780
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3058 5488 3538
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5828 3058 5856 3334
rect 5920 3194 5948 4014
rect 6012 3602 6040 4150
rect 6748 4146 7420 4162
rect 6748 4140 7432 4146
rect 6748 4134 7380 4140
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6104 3670 6132 4014
rect 6472 3913 6500 4014
rect 6644 3936 6696 3942
rect 6458 3904 6514 3913
rect 6644 3878 6696 3884
rect 6458 3839 6514 3848
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6012 3058 6040 3538
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6104 3126 6132 3470
rect 6198 3292 6506 3301
rect 6198 3290 6204 3292
rect 6260 3290 6284 3292
rect 6340 3290 6364 3292
rect 6420 3290 6444 3292
rect 6500 3290 6506 3292
rect 6260 3238 6262 3290
rect 6442 3238 6444 3290
rect 6198 3236 6204 3238
rect 6260 3236 6284 3238
rect 6340 3236 6364 3238
rect 6420 3236 6444 3238
rect 6500 3236 6506 3238
rect 6198 3227 6506 3236
rect 6656 3194 6684 3878
rect 6748 3534 6776 4134
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6840 3738 6868 4014
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3670 6960 3878
rect 7116 3738 7144 3946
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 6920 3664 6972 3670
rect 7208 3618 7236 3946
rect 6920 3606 6972 3612
rect 7116 3602 7236 3618
rect 7300 3602 7328 4134
rect 7380 4082 7432 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7576 3942 7604 4082
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7760 3602 7788 4082
rect 8036 3738 8064 4082
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7104 3596 7236 3602
rect 7156 3590 7236 3596
rect 7288 3596 7340 3602
rect 7104 3538 7156 3544
rect 7288 3538 7340 3544
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 6736 3528 6788 3534
rect 7196 3528 7248 3534
rect 6736 3470 6788 3476
rect 7194 3496 7196 3505
rect 7248 3496 7250 3505
rect 6920 3460 6972 3466
rect 7194 3431 7250 3440
rect 6920 3402 6972 3408
rect 6932 3194 6960 3402
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 5224 3012 5304 3040
rect 5356 3052 5408 3058
rect 5172 2994 5224 3000
rect 5356 2994 5408 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5184 2650 5212 2790
rect 5538 2748 5846 2757
rect 5538 2746 5544 2748
rect 5600 2746 5624 2748
rect 5680 2746 5704 2748
rect 5760 2746 5784 2748
rect 5840 2746 5846 2748
rect 5600 2694 5602 2746
rect 5782 2694 5784 2746
rect 5538 2692 5544 2694
rect 5600 2692 5624 2694
rect 5680 2692 5704 2694
rect 5760 2692 5784 2694
rect 5840 2692 5846 2694
rect 5538 2683 5846 2692
rect 6012 2650 6040 2994
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6104 2446 6132 3062
rect 7484 3058 7512 3334
rect 7760 3194 7788 3538
rect 8128 3194 8156 4082
rect 8220 3534 8248 4966
rect 8312 3913 8340 5102
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8404 3942 8432 4082
rect 8496 3942 8524 5170
rect 8597 4924 8905 4933
rect 8597 4922 8603 4924
rect 8659 4922 8683 4924
rect 8739 4922 8763 4924
rect 8819 4922 8843 4924
rect 8899 4922 8905 4924
rect 8659 4870 8661 4922
rect 8841 4870 8843 4922
rect 8597 4868 8603 4870
rect 8659 4868 8683 4870
rect 8739 4868 8763 4870
rect 8819 4868 8843 4870
rect 8899 4868 8905 4870
rect 8597 4859 8905 4868
rect 9232 4826 9260 5170
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9257 4380 9565 4389
rect 9257 4378 9263 4380
rect 9319 4378 9343 4380
rect 9399 4378 9423 4380
rect 9479 4378 9503 4380
rect 9559 4378 9565 4380
rect 9319 4326 9321 4378
rect 9501 4326 9503 4378
rect 9257 4324 9263 4326
rect 9319 4324 9343 4326
rect 9399 4324 9423 4326
rect 9479 4324 9503 4326
rect 9559 4324 9565 4326
rect 9257 4315 9565 4324
rect 9784 4146 9812 4966
rect 9876 4146 9904 5102
rect 10704 4622 10732 5238
rect 10980 5222 11100 5238
rect 10980 5114 11008 5222
rect 10888 5086 11008 5114
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10888 4282 10916 5086
rect 11164 4622 11192 6734
rect 11440 5166 11468 7278
rect 11656 7100 11964 7109
rect 11656 7098 11662 7100
rect 11718 7098 11742 7100
rect 11798 7098 11822 7100
rect 11878 7098 11902 7100
rect 11958 7098 11964 7100
rect 11718 7046 11720 7098
rect 11900 7046 11902 7098
rect 11656 7044 11662 7046
rect 11718 7044 11742 7046
rect 11798 7044 11822 7046
rect 11878 7044 11902 7046
rect 11958 7044 11964 7046
rect 11656 7035 11964 7044
rect 11992 6322 12020 9522
rect 12176 9178 12204 10118
rect 12360 9926 12388 10610
rect 12636 10062 12664 10678
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10169 13032 10542
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12316 9820 12624 9829
rect 12316 9818 12322 9820
rect 12378 9818 12402 9820
rect 12458 9818 12482 9820
rect 12538 9818 12562 9820
rect 12618 9818 12624 9820
rect 12378 9766 12380 9818
rect 12560 9766 12562 9818
rect 12316 9764 12322 9766
rect 12378 9764 12402 9766
rect 12458 9764 12482 9766
rect 12538 9764 12562 9766
rect 12618 9764 12624 9766
rect 12316 9755 12624 9764
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8634 12204 8910
rect 12316 8732 12624 8741
rect 12316 8730 12322 8732
rect 12378 8730 12402 8732
rect 12458 8730 12482 8732
rect 12538 8730 12562 8732
rect 12618 8730 12624 8732
rect 12378 8678 12380 8730
rect 12560 8678 12562 8730
rect 12316 8676 12322 8678
rect 12378 8676 12402 8678
rect 12458 8676 12482 8678
rect 12538 8676 12562 8678
rect 12618 8676 12624 8678
rect 12316 8667 12624 8676
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12084 7410 12112 8434
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7818 12480 8230
rect 12912 8090 12940 8366
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12316 7644 12624 7653
rect 12316 7642 12322 7644
rect 12378 7642 12402 7644
rect 12458 7642 12482 7644
rect 12538 7642 12562 7644
rect 12618 7642 12624 7644
rect 12378 7590 12380 7642
rect 12560 7590 12562 7642
rect 12316 7588 12322 7590
rect 12378 7588 12402 7590
rect 12458 7588 12482 7590
rect 12538 7588 12562 7590
rect 12618 7588 12624 7590
rect 12316 7579 12624 7588
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6730 12480 7142
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12316 6556 12624 6565
rect 12316 6554 12322 6556
rect 12378 6554 12402 6556
rect 12458 6554 12482 6556
rect 12538 6554 12562 6556
rect 12618 6554 12624 6556
rect 12378 6502 12380 6554
rect 12560 6502 12562 6554
rect 12316 6500 12322 6502
rect 12378 6500 12402 6502
rect 12458 6500 12482 6502
rect 12538 6500 12562 6502
rect 12618 6500 12624 6502
rect 12316 6491 12624 6500
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 6089 13032 6190
rect 12990 6080 13046 6089
rect 11656 6012 11964 6021
rect 12990 6015 13046 6024
rect 11656 6010 11662 6012
rect 11718 6010 11742 6012
rect 11798 6010 11822 6012
rect 11878 6010 11902 6012
rect 11958 6010 11964 6012
rect 11718 5958 11720 6010
rect 11900 5958 11902 6010
rect 11656 5956 11662 5958
rect 11718 5956 11742 5958
rect 11798 5956 11822 5958
rect 11878 5956 11902 5958
rect 11958 5956 11964 5958
rect 11656 5947 11964 5956
rect 12316 5468 12624 5477
rect 12316 5466 12322 5468
rect 12378 5466 12402 5468
rect 12458 5466 12482 5468
rect 12538 5466 12562 5468
rect 12618 5466 12624 5468
rect 12378 5414 12380 5466
rect 12560 5414 12562 5466
rect 12316 5412 12322 5414
rect 12378 5412 12402 5414
rect 12458 5412 12482 5414
rect 12538 5412 12562 5414
rect 12618 5412 12624 5414
rect 12316 5403 12624 5412
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10980 4282 11008 4490
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 8392 3936 8444 3942
rect 8298 3904 8354 3913
rect 8392 3878 8444 3884
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8298 3839 8354 3848
rect 8404 3720 8432 3878
rect 8597 3836 8905 3845
rect 8597 3834 8603 3836
rect 8659 3834 8683 3836
rect 8739 3834 8763 3836
rect 8819 3834 8843 3836
rect 8899 3834 8905 3836
rect 8659 3782 8661 3834
rect 8841 3782 8843 3834
rect 8597 3780 8603 3782
rect 8659 3780 8683 3782
rect 8739 3780 8763 3782
rect 8819 3780 8843 3782
rect 8899 3780 8905 3782
rect 8597 3771 8905 3780
rect 8404 3692 8892 3720
rect 8864 3602 8892 3692
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8208 3528 8260 3534
rect 8392 3528 8444 3534
rect 8208 3470 8260 3476
rect 8298 3496 8354 3505
rect 8354 3476 8392 3482
rect 8354 3470 8444 3476
rect 8354 3454 8432 3470
rect 8298 3431 8354 3440
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8220 3194 8248 3334
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8312 3058 8340 3334
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 6472 2650 6500 2994
rect 8404 2922 8432 3454
rect 8496 3058 8524 3538
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8588 3194 8616 3470
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8484 3052 8536 3058
rect 8680 3040 8708 3470
rect 8956 3466 8984 3878
rect 9048 3534 9076 3878
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3074 9076 3334
rect 9140 3194 9168 3946
rect 9232 3738 9260 3946
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9784 3670 9812 4082
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3398 9352 3470
rect 9416 3398 9444 3606
rect 9600 3534 9628 3606
rect 9784 3534 9812 3606
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9257 3292 9565 3301
rect 9257 3290 9263 3292
rect 9319 3290 9343 3292
rect 9399 3290 9423 3292
rect 9479 3290 9503 3292
rect 9559 3290 9565 3292
rect 9319 3238 9321 3290
rect 9501 3238 9503 3290
rect 9257 3236 9263 3238
rect 9319 3236 9343 3238
rect 9399 3236 9423 3238
rect 9479 3236 9503 3238
rect 9559 3236 9565 3238
rect 9257 3227 9565 3236
rect 9692 3194 9720 3470
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9312 3120 9364 3126
rect 9048 3068 9312 3074
rect 9048 3062 9364 3068
rect 8536 3012 8708 3040
rect 8944 3052 8996 3058
rect 8484 2994 8536 3000
rect 9048 3046 9352 3062
rect 9784 3058 9812 3470
rect 10428 3126 10456 3946
rect 10704 3738 10732 4014
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10796 3618 10824 3878
rect 10888 3738 10916 4082
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10796 3590 10916 3618
rect 10888 3534 10916 3590
rect 10980 3534 11008 4218
rect 11072 4214 11100 4422
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11164 3602 11192 4558
rect 11256 4078 11284 4966
rect 11440 4826 11468 5102
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11532 4690 11560 4966
rect 11656 4924 11964 4933
rect 11656 4922 11662 4924
rect 11718 4922 11742 4924
rect 11798 4922 11822 4924
rect 11878 4922 11902 4924
rect 11958 4922 11964 4924
rect 11718 4870 11720 4922
rect 11900 4870 11902 4922
rect 11656 4868 11662 4870
rect 11718 4868 11742 4870
rect 11798 4868 11822 4870
rect 11878 4868 11902 4870
rect 11958 4868 11964 4870
rect 11656 4859 11964 4868
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 12176 4554 12204 4966
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11348 4282 11376 4422
rect 12316 4380 12624 4389
rect 12316 4378 12322 4380
rect 12378 4378 12402 4380
rect 12458 4378 12482 4380
rect 12538 4378 12562 4380
rect 12618 4378 12624 4380
rect 12378 4326 12380 4378
rect 12560 4326 12562 4378
rect 12316 4324 12322 4326
rect 12378 4324 12402 4326
rect 12458 4324 12482 4326
rect 12538 4324 12562 4326
rect 12618 4324 12624 4326
rect 12316 4315 12624 4324
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11656 3836 11964 3845
rect 11656 3834 11662 3836
rect 11718 3834 11742 3836
rect 11798 3834 11822 3836
rect 11878 3834 11902 3836
rect 11958 3834 11964 3836
rect 11718 3782 11720 3834
rect 11900 3782 11902 3834
rect 11656 3780 11662 3782
rect 11718 3780 11742 3782
rect 11798 3780 11822 3782
rect 11878 3780 11902 3782
rect 11958 3780 11964 3782
rect 11656 3771 11964 3780
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 9772 3052 9824 3058
rect 8944 2994 8996 3000
rect 9772 2994 9824 3000
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8597 2748 8905 2757
rect 8597 2746 8603 2748
rect 8659 2746 8683 2748
rect 8739 2746 8763 2748
rect 8819 2746 8843 2748
rect 8899 2746 8905 2748
rect 8659 2694 8661 2746
rect 8841 2694 8843 2746
rect 8597 2692 8603 2694
rect 8659 2692 8683 2694
rect 8739 2692 8763 2694
rect 8819 2692 8843 2694
rect 8899 2692 8905 2694
rect 8597 2683 8905 2692
rect 8956 2650 8984 2994
rect 10888 2990 10916 3470
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10428 2650 10456 2926
rect 11072 2922 11100 3334
rect 12084 3058 12112 3878
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 3194 12204 3334
rect 12316 3292 12624 3301
rect 12316 3290 12322 3292
rect 12378 3290 12402 3292
rect 12458 3290 12482 3292
rect 12538 3290 12562 3292
rect 12618 3290 12624 3292
rect 12378 3238 12380 3290
rect 12560 3238 12562 3290
rect 12316 3236 12322 3238
rect 12378 3236 12402 3238
rect 12458 3236 12482 3238
rect 12538 3236 12562 3238
rect 12618 3236 12624 3238
rect 12316 3227 12624 3236
rect 12728 3194 12756 3402
rect 12820 3194 12848 4762
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3738 12940 4082
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 11072 2514 11100 2858
rect 11656 2748 11964 2757
rect 11656 2746 11662 2748
rect 11718 2746 11742 2748
rect 11798 2746 11822 2748
rect 11878 2746 11902 2748
rect 11958 2746 11964 2748
rect 11718 2694 11720 2746
rect 11900 2694 11902 2746
rect 11656 2692 11662 2694
rect 11718 2692 11742 2694
rect 11798 2692 11822 2694
rect 11878 2692 11902 2694
rect 11958 2692 11964 2694
rect 11656 2683 11964 2692
rect 13096 2650 13124 9318
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 940 2440 992 2446
rect 2596 2440 2648 2446
rect 940 2382 992 2388
rect 2516 2400 2596 2428
rect 952 800 980 2382
rect 2516 800 2544 2400
rect 4160 2440 4212 2446
rect 2596 2382 2648 2388
rect 4080 2400 4160 2428
rect 3139 2204 3447 2213
rect 3139 2202 3145 2204
rect 3201 2202 3225 2204
rect 3281 2202 3305 2204
rect 3361 2202 3385 2204
rect 3441 2202 3447 2204
rect 3201 2150 3203 2202
rect 3383 2150 3385 2202
rect 3139 2148 3145 2150
rect 3201 2148 3225 2150
rect 3281 2148 3305 2150
rect 3361 2148 3385 2150
rect 3441 2148 3447 2150
rect 3139 2139 3447 2148
rect 4080 800 4108 2400
rect 5724 2440 5776 2446
rect 4160 2382 4212 2388
rect 5644 2400 5724 2428
rect 5644 800 5672 2400
rect 5724 2382 5776 2388
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 6198 2204 6506 2213
rect 6198 2202 6204 2204
rect 6260 2202 6284 2204
rect 6340 2202 6364 2204
rect 6420 2202 6444 2204
rect 6500 2202 6506 2204
rect 6260 2150 6262 2202
rect 6442 2150 6444 2202
rect 6198 2148 6204 2150
rect 6260 2148 6284 2150
rect 6340 2148 6364 2150
rect 6420 2148 6444 2150
rect 6500 2148 6506 2150
rect 6198 2139 6506 2148
rect 7208 800 7236 2382
rect 8772 800 8800 2382
rect 9257 2204 9565 2213
rect 9257 2202 9263 2204
rect 9319 2202 9343 2204
rect 9399 2202 9423 2204
rect 9479 2202 9503 2204
rect 9559 2202 9565 2204
rect 9319 2150 9321 2202
rect 9501 2150 9503 2202
rect 9257 2148 9263 2150
rect 9319 2148 9343 2150
rect 9399 2148 9423 2150
rect 9479 2148 9503 2150
rect 9559 2148 9565 2150
rect 9257 2139 9565 2148
rect 10336 800 10364 2382
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 11900 800 11928 2314
rect 12316 2204 12624 2213
rect 12316 2202 12322 2204
rect 12378 2202 12402 2204
rect 12458 2202 12482 2204
rect 12538 2202 12562 2204
rect 12618 2202 12624 2204
rect 12378 2150 12380 2202
rect 12560 2150 12562 2202
rect 12316 2148 12322 2150
rect 12378 2148 12402 2150
rect 12458 2148 12482 2150
rect 12538 2148 12562 2150
rect 12618 2148 12624 2150
rect 12316 2139 12624 2148
rect 13280 2009 13308 2314
rect 13266 2000 13322 2009
rect 13266 1935 13322 1944
rect 13464 800 13492 2994
rect 938 0 994 800
rect 2502 0 2558 800
rect 4066 0 4122 800
rect 5630 0 5686 800
rect 7194 0 7250 800
rect 8758 0 8814 800
rect 10322 0 10378 800
rect 11886 0 11942 800
rect 13450 0 13506 800
<< via2 >>
rect 3145 14170 3201 14172
rect 3225 14170 3281 14172
rect 3305 14170 3361 14172
rect 3385 14170 3441 14172
rect 3145 14118 3191 14170
rect 3191 14118 3201 14170
rect 3225 14118 3255 14170
rect 3255 14118 3267 14170
rect 3267 14118 3281 14170
rect 3305 14118 3319 14170
rect 3319 14118 3331 14170
rect 3331 14118 3361 14170
rect 3385 14118 3395 14170
rect 3395 14118 3441 14170
rect 3145 14116 3201 14118
rect 3225 14116 3281 14118
rect 3305 14116 3361 14118
rect 3385 14116 3441 14118
rect 6204 14170 6260 14172
rect 6284 14170 6340 14172
rect 6364 14170 6420 14172
rect 6444 14170 6500 14172
rect 6204 14118 6250 14170
rect 6250 14118 6260 14170
rect 6284 14118 6314 14170
rect 6314 14118 6326 14170
rect 6326 14118 6340 14170
rect 6364 14118 6378 14170
rect 6378 14118 6390 14170
rect 6390 14118 6420 14170
rect 6444 14118 6454 14170
rect 6454 14118 6500 14170
rect 6204 14116 6260 14118
rect 6284 14116 6340 14118
rect 6364 14116 6420 14118
rect 6444 14116 6500 14118
rect 9263 14170 9319 14172
rect 9343 14170 9399 14172
rect 9423 14170 9479 14172
rect 9503 14170 9559 14172
rect 9263 14118 9309 14170
rect 9309 14118 9319 14170
rect 9343 14118 9373 14170
rect 9373 14118 9385 14170
rect 9385 14118 9399 14170
rect 9423 14118 9437 14170
rect 9437 14118 9449 14170
rect 9449 14118 9479 14170
rect 9503 14118 9513 14170
rect 9513 14118 9559 14170
rect 9263 14116 9319 14118
rect 9343 14116 9399 14118
rect 9423 14116 9479 14118
rect 9503 14116 9559 14118
rect 13266 14184 13322 14240
rect 12322 14170 12378 14172
rect 12402 14170 12458 14172
rect 12482 14170 12538 14172
rect 12562 14170 12618 14172
rect 12322 14118 12368 14170
rect 12368 14118 12378 14170
rect 12402 14118 12432 14170
rect 12432 14118 12444 14170
rect 12444 14118 12458 14170
rect 12482 14118 12496 14170
rect 12496 14118 12508 14170
rect 12508 14118 12538 14170
rect 12562 14118 12572 14170
rect 12572 14118 12618 14170
rect 12322 14116 12378 14118
rect 12402 14116 12458 14118
rect 12482 14116 12538 14118
rect 12562 14116 12618 14118
rect 2485 13626 2541 13628
rect 2565 13626 2621 13628
rect 2645 13626 2701 13628
rect 2725 13626 2781 13628
rect 2485 13574 2531 13626
rect 2531 13574 2541 13626
rect 2565 13574 2595 13626
rect 2595 13574 2607 13626
rect 2607 13574 2621 13626
rect 2645 13574 2659 13626
rect 2659 13574 2671 13626
rect 2671 13574 2701 13626
rect 2725 13574 2735 13626
rect 2735 13574 2781 13626
rect 2485 13572 2541 13574
rect 2565 13572 2621 13574
rect 2645 13572 2701 13574
rect 2725 13572 2781 13574
rect 3145 13082 3201 13084
rect 3225 13082 3281 13084
rect 3305 13082 3361 13084
rect 3385 13082 3441 13084
rect 3145 13030 3191 13082
rect 3191 13030 3201 13082
rect 3225 13030 3255 13082
rect 3255 13030 3267 13082
rect 3267 13030 3281 13082
rect 3305 13030 3319 13082
rect 3319 13030 3331 13082
rect 3331 13030 3361 13082
rect 3385 13030 3395 13082
rect 3395 13030 3441 13082
rect 3145 13028 3201 13030
rect 3225 13028 3281 13030
rect 3305 13028 3361 13030
rect 3385 13028 3441 13030
rect 2485 12538 2541 12540
rect 2565 12538 2621 12540
rect 2645 12538 2701 12540
rect 2725 12538 2781 12540
rect 2485 12486 2531 12538
rect 2531 12486 2541 12538
rect 2565 12486 2595 12538
rect 2595 12486 2607 12538
rect 2607 12486 2621 12538
rect 2645 12486 2659 12538
rect 2659 12486 2671 12538
rect 2671 12486 2701 12538
rect 2725 12486 2735 12538
rect 2735 12486 2781 12538
rect 2485 12484 2541 12486
rect 2565 12484 2621 12486
rect 2645 12484 2701 12486
rect 2725 12484 2781 12486
rect 4066 12280 4122 12336
rect 3145 11994 3201 11996
rect 3225 11994 3281 11996
rect 3305 11994 3361 11996
rect 3385 11994 3441 11996
rect 3145 11942 3191 11994
rect 3191 11942 3201 11994
rect 3225 11942 3255 11994
rect 3255 11942 3267 11994
rect 3267 11942 3281 11994
rect 3305 11942 3319 11994
rect 3319 11942 3331 11994
rect 3331 11942 3361 11994
rect 3385 11942 3395 11994
rect 3395 11942 3441 11994
rect 3145 11940 3201 11942
rect 3225 11940 3281 11942
rect 3305 11940 3361 11942
rect 3385 11940 3441 11942
rect 2485 11450 2541 11452
rect 2565 11450 2621 11452
rect 2645 11450 2701 11452
rect 2725 11450 2781 11452
rect 2485 11398 2531 11450
rect 2531 11398 2541 11450
rect 2565 11398 2595 11450
rect 2595 11398 2607 11450
rect 2607 11398 2621 11450
rect 2645 11398 2659 11450
rect 2659 11398 2671 11450
rect 2671 11398 2701 11450
rect 2725 11398 2735 11450
rect 2735 11398 2781 11450
rect 2485 11396 2541 11398
rect 2565 11396 2621 11398
rect 2645 11396 2701 11398
rect 2725 11396 2781 11398
rect 3145 10906 3201 10908
rect 3225 10906 3281 10908
rect 3305 10906 3361 10908
rect 3385 10906 3441 10908
rect 3145 10854 3191 10906
rect 3191 10854 3201 10906
rect 3225 10854 3255 10906
rect 3255 10854 3267 10906
rect 3267 10854 3281 10906
rect 3305 10854 3319 10906
rect 3319 10854 3331 10906
rect 3331 10854 3361 10906
rect 3385 10854 3395 10906
rect 3395 10854 3441 10906
rect 3145 10852 3201 10854
rect 3225 10852 3281 10854
rect 3305 10852 3361 10854
rect 3385 10852 3441 10854
rect 2485 10362 2541 10364
rect 2565 10362 2621 10364
rect 2645 10362 2701 10364
rect 2725 10362 2781 10364
rect 2485 10310 2531 10362
rect 2531 10310 2541 10362
rect 2565 10310 2595 10362
rect 2595 10310 2607 10362
rect 2607 10310 2621 10362
rect 2645 10310 2659 10362
rect 2659 10310 2671 10362
rect 2671 10310 2701 10362
rect 2725 10310 2735 10362
rect 2735 10310 2781 10362
rect 2485 10308 2541 10310
rect 2565 10308 2621 10310
rect 2645 10308 2701 10310
rect 2725 10308 2781 10310
rect 3145 9818 3201 9820
rect 3225 9818 3281 9820
rect 3305 9818 3361 9820
rect 3385 9818 3441 9820
rect 3145 9766 3191 9818
rect 3191 9766 3201 9818
rect 3225 9766 3255 9818
rect 3255 9766 3267 9818
rect 3267 9766 3281 9818
rect 3305 9766 3319 9818
rect 3319 9766 3331 9818
rect 3331 9766 3361 9818
rect 3385 9766 3395 9818
rect 3395 9766 3441 9818
rect 3145 9764 3201 9766
rect 3225 9764 3281 9766
rect 3305 9764 3361 9766
rect 3385 9764 3441 9766
rect 2485 9274 2541 9276
rect 2565 9274 2621 9276
rect 2645 9274 2701 9276
rect 2725 9274 2781 9276
rect 2485 9222 2531 9274
rect 2531 9222 2541 9274
rect 2565 9222 2595 9274
rect 2595 9222 2607 9274
rect 2607 9222 2621 9274
rect 2645 9222 2659 9274
rect 2659 9222 2671 9274
rect 2671 9222 2701 9274
rect 2725 9222 2735 9274
rect 2735 9222 2781 9274
rect 2485 9220 2541 9222
rect 2565 9220 2621 9222
rect 2645 9220 2701 9222
rect 2725 9220 2781 9222
rect 3145 8730 3201 8732
rect 3225 8730 3281 8732
rect 3305 8730 3361 8732
rect 3385 8730 3441 8732
rect 3145 8678 3191 8730
rect 3191 8678 3201 8730
rect 3225 8678 3255 8730
rect 3255 8678 3267 8730
rect 3267 8678 3281 8730
rect 3305 8678 3319 8730
rect 3319 8678 3331 8730
rect 3331 8678 3361 8730
rect 3385 8678 3395 8730
rect 3395 8678 3441 8730
rect 3145 8676 3201 8678
rect 3225 8676 3281 8678
rect 3305 8676 3361 8678
rect 3385 8676 3441 8678
rect 938 4120 994 4176
rect 2485 8186 2541 8188
rect 2565 8186 2621 8188
rect 2645 8186 2701 8188
rect 2725 8186 2781 8188
rect 2485 8134 2531 8186
rect 2531 8134 2541 8186
rect 2565 8134 2595 8186
rect 2595 8134 2607 8186
rect 2607 8134 2621 8186
rect 2645 8134 2659 8186
rect 2659 8134 2671 8186
rect 2671 8134 2701 8186
rect 2725 8134 2735 8186
rect 2735 8134 2781 8186
rect 2485 8132 2541 8134
rect 2565 8132 2621 8134
rect 2645 8132 2701 8134
rect 2725 8132 2781 8134
rect 3145 7642 3201 7644
rect 3225 7642 3281 7644
rect 3305 7642 3361 7644
rect 3385 7642 3441 7644
rect 3145 7590 3191 7642
rect 3191 7590 3201 7642
rect 3225 7590 3255 7642
rect 3255 7590 3267 7642
rect 3267 7590 3281 7642
rect 3305 7590 3319 7642
rect 3319 7590 3331 7642
rect 3331 7590 3361 7642
rect 3385 7590 3395 7642
rect 3395 7590 3441 7642
rect 3145 7588 3201 7590
rect 3225 7588 3281 7590
rect 3305 7588 3361 7590
rect 3385 7588 3441 7590
rect 2485 7098 2541 7100
rect 2565 7098 2621 7100
rect 2645 7098 2701 7100
rect 2725 7098 2781 7100
rect 2485 7046 2531 7098
rect 2531 7046 2541 7098
rect 2565 7046 2595 7098
rect 2595 7046 2607 7098
rect 2607 7046 2621 7098
rect 2645 7046 2659 7098
rect 2659 7046 2671 7098
rect 2671 7046 2701 7098
rect 2725 7046 2735 7098
rect 2735 7046 2781 7098
rect 2485 7044 2541 7046
rect 2565 7044 2621 7046
rect 2645 7044 2701 7046
rect 2725 7044 2781 7046
rect 2485 6010 2541 6012
rect 2565 6010 2621 6012
rect 2645 6010 2701 6012
rect 2725 6010 2781 6012
rect 2485 5958 2531 6010
rect 2531 5958 2541 6010
rect 2565 5958 2595 6010
rect 2595 5958 2607 6010
rect 2607 5958 2621 6010
rect 2645 5958 2659 6010
rect 2659 5958 2671 6010
rect 2671 5958 2701 6010
rect 2725 5958 2735 6010
rect 2735 5958 2781 6010
rect 2485 5956 2541 5958
rect 2565 5956 2621 5958
rect 2645 5956 2701 5958
rect 2725 5956 2781 5958
rect 2485 4922 2541 4924
rect 2565 4922 2621 4924
rect 2645 4922 2701 4924
rect 2725 4922 2781 4924
rect 2485 4870 2531 4922
rect 2531 4870 2541 4922
rect 2565 4870 2595 4922
rect 2595 4870 2607 4922
rect 2607 4870 2621 4922
rect 2645 4870 2659 4922
rect 2659 4870 2671 4922
rect 2671 4870 2701 4922
rect 2725 4870 2735 4922
rect 2735 4870 2781 4922
rect 2485 4868 2541 4870
rect 2565 4868 2621 4870
rect 2645 4868 2701 4870
rect 2725 4868 2781 4870
rect 2686 4020 2688 4040
rect 2688 4020 2740 4040
rect 2740 4020 2742 4040
rect 2686 3984 2742 4020
rect 3145 6554 3201 6556
rect 3225 6554 3281 6556
rect 3305 6554 3361 6556
rect 3385 6554 3441 6556
rect 3145 6502 3191 6554
rect 3191 6502 3201 6554
rect 3225 6502 3255 6554
rect 3255 6502 3267 6554
rect 3267 6502 3281 6554
rect 3305 6502 3319 6554
rect 3319 6502 3331 6554
rect 3331 6502 3361 6554
rect 3385 6502 3395 6554
rect 3395 6502 3441 6554
rect 3145 6500 3201 6502
rect 3225 6500 3281 6502
rect 3305 6500 3361 6502
rect 3385 6500 3441 6502
rect 3145 5466 3201 5468
rect 3225 5466 3281 5468
rect 3305 5466 3361 5468
rect 3385 5466 3441 5468
rect 3145 5414 3191 5466
rect 3191 5414 3201 5466
rect 3225 5414 3255 5466
rect 3255 5414 3267 5466
rect 3267 5414 3281 5466
rect 3305 5414 3319 5466
rect 3319 5414 3331 5466
rect 3331 5414 3361 5466
rect 3385 5414 3395 5466
rect 3395 5414 3441 5466
rect 3145 5412 3201 5414
rect 3225 5412 3281 5414
rect 3305 5412 3361 5414
rect 3385 5412 3441 5414
rect 3145 4378 3201 4380
rect 3225 4378 3281 4380
rect 3305 4378 3361 4380
rect 3385 4378 3441 4380
rect 3145 4326 3191 4378
rect 3191 4326 3201 4378
rect 3225 4326 3255 4378
rect 3255 4326 3267 4378
rect 3267 4326 3281 4378
rect 3305 4326 3319 4378
rect 3319 4326 3331 4378
rect 3331 4326 3361 4378
rect 3385 4326 3395 4378
rect 3395 4326 3441 4378
rect 3145 4324 3201 4326
rect 3225 4324 3281 4326
rect 3305 4324 3361 4326
rect 3385 4324 3441 4326
rect 2485 3834 2541 3836
rect 2565 3834 2621 3836
rect 2645 3834 2701 3836
rect 2725 3834 2781 3836
rect 2485 3782 2531 3834
rect 2531 3782 2541 3834
rect 2565 3782 2595 3834
rect 2595 3782 2607 3834
rect 2607 3782 2621 3834
rect 2645 3782 2659 3834
rect 2659 3782 2671 3834
rect 2671 3782 2701 3834
rect 2725 3782 2735 3834
rect 2735 3782 2781 3834
rect 2485 3780 2541 3782
rect 2565 3780 2621 3782
rect 2645 3780 2701 3782
rect 2725 3780 2781 3782
rect 3145 3290 3201 3292
rect 3225 3290 3281 3292
rect 3305 3290 3361 3292
rect 3385 3290 3441 3292
rect 3145 3238 3191 3290
rect 3191 3238 3201 3290
rect 3225 3238 3255 3290
rect 3255 3238 3267 3290
rect 3267 3238 3281 3290
rect 3305 3238 3319 3290
rect 3319 3238 3331 3290
rect 3331 3238 3361 3290
rect 3385 3238 3395 3290
rect 3395 3238 3441 3290
rect 3145 3236 3201 3238
rect 3225 3236 3281 3238
rect 3305 3236 3361 3238
rect 3385 3236 3441 3238
rect 2485 2746 2541 2748
rect 2565 2746 2621 2748
rect 2645 2746 2701 2748
rect 2725 2746 2781 2748
rect 2485 2694 2531 2746
rect 2531 2694 2541 2746
rect 2565 2694 2595 2746
rect 2595 2694 2607 2746
rect 2607 2694 2621 2746
rect 2645 2694 2659 2746
rect 2659 2694 2671 2746
rect 2671 2694 2701 2746
rect 2725 2694 2735 2746
rect 2735 2694 2781 2746
rect 2485 2692 2541 2694
rect 2565 2692 2621 2694
rect 2645 2692 2701 2694
rect 2725 2692 2781 2694
rect 5544 13626 5600 13628
rect 5624 13626 5680 13628
rect 5704 13626 5760 13628
rect 5784 13626 5840 13628
rect 5544 13574 5590 13626
rect 5590 13574 5600 13626
rect 5624 13574 5654 13626
rect 5654 13574 5666 13626
rect 5666 13574 5680 13626
rect 5704 13574 5718 13626
rect 5718 13574 5730 13626
rect 5730 13574 5760 13626
rect 5784 13574 5794 13626
rect 5794 13574 5840 13626
rect 5544 13572 5600 13574
rect 5624 13572 5680 13574
rect 5704 13572 5760 13574
rect 5784 13572 5840 13574
rect 8603 13626 8659 13628
rect 8683 13626 8739 13628
rect 8763 13626 8819 13628
rect 8843 13626 8899 13628
rect 8603 13574 8649 13626
rect 8649 13574 8659 13626
rect 8683 13574 8713 13626
rect 8713 13574 8725 13626
rect 8725 13574 8739 13626
rect 8763 13574 8777 13626
rect 8777 13574 8789 13626
rect 8789 13574 8819 13626
rect 8843 13574 8853 13626
rect 8853 13574 8899 13626
rect 8603 13572 8659 13574
rect 8683 13572 8739 13574
rect 8763 13572 8819 13574
rect 8843 13572 8899 13574
rect 6204 13082 6260 13084
rect 6284 13082 6340 13084
rect 6364 13082 6420 13084
rect 6444 13082 6500 13084
rect 6204 13030 6250 13082
rect 6250 13030 6260 13082
rect 6284 13030 6314 13082
rect 6314 13030 6326 13082
rect 6326 13030 6340 13082
rect 6364 13030 6378 13082
rect 6378 13030 6390 13082
rect 6390 13030 6420 13082
rect 6444 13030 6454 13082
rect 6454 13030 6500 13082
rect 6204 13028 6260 13030
rect 6284 13028 6340 13030
rect 6364 13028 6420 13030
rect 6444 13028 6500 13030
rect 5544 12538 5600 12540
rect 5624 12538 5680 12540
rect 5704 12538 5760 12540
rect 5784 12538 5840 12540
rect 5544 12486 5590 12538
rect 5590 12486 5600 12538
rect 5624 12486 5654 12538
rect 5654 12486 5666 12538
rect 5666 12486 5680 12538
rect 5704 12486 5718 12538
rect 5718 12486 5730 12538
rect 5730 12486 5760 12538
rect 5784 12486 5794 12538
rect 5794 12486 5840 12538
rect 5544 12484 5600 12486
rect 5624 12484 5680 12486
rect 5704 12484 5760 12486
rect 5784 12484 5840 12486
rect 6204 11994 6260 11996
rect 6284 11994 6340 11996
rect 6364 11994 6420 11996
rect 6444 11994 6500 11996
rect 6204 11942 6250 11994
rect 6250 11942 6260 11994
rect 6284 11942 6314 11994
rect 6314 11942 6326 11994
rect 6326 11942 6340 11994
rect 6364 11942 6378 11994
rect 6378 11942 6390 11994
rect 6390 11942 6420 11994
rect 6444 11942 6454 11994
rect 6454 11942 6500 11994
rect 6204 11940 6260 11942
rect 6284 11940 6340 11942
rect 6364 11940 6420 11942
rect 6444 11940 6500 11942
rect 5544 11450 5600 11452
rect 5624 11450 5680 11452
rect 5704 11450 5760 11452
rect 5784 11450 5840 11452
rect 5544 11398 5590 11450
rect 5590 11398 5600 11450
rect 5624 11398 5654 11450
rect 5654 11398 5666 11450
rect 5666 11398 5680 11450
rect 5704 11398 5718 11450
rect 5718 11398 5730 11450
rect 5730 11398 5760 11450
rect 5784 11398 5794 11450
rect 5794 11398 5840 11450
rect 5544 11396 5600 11398
rect 5624 11396 5680 11398
rect 5704 11396 5760 11398
rect 5784 11396 5840 11398
rect 5544 10362 5600 10364
rect 5624 10362 5680 10364
rect 5704 10362 5760 10364
rect 5784 10362 5840 10364
rect 5544 10310 5590 10362
rect 5590 10310 5600 10362
rect 5624 10310 5654 10362
rect 5654 10310 5666 10362
rect 5666 10310 5680 10362
rect 5704 10310 5718 10362
rect 5718 10310 5730 10362
rect 5730 10310 5760 10362
rect 5784 10310 5794 10362
rect 5794 10310 5840 10362
rect 5544 10308 5600 10310
rect 5624 10308 5680 10310
rect 5704 10308 5760 10310
rect 5784 10308 5840 10310
rect 5544 9274 5600 9276
rect 5624 9274 5680 9276
rect 5704 9274 5760 9276
rect 5784 9274 5840 9276
rect 5544 9222 5590 9274
rect 5590 9222 5600 9274
rect 5624 9222 5654 9274
rect 5654 9222 5666 9274
rect 5666 9222 5680 9274
rect 5704 9222 5718 9274
rect 5718 9222 5730 9274
rect 5730 9222 5760 9274
rect 5784 9222 5794 9274
rect 5794 9222 5840 9274
rect 5544 9220 5600 9222
rect 5624 9220 5680 9222
rect 5704 9220 5760 9222
rect 5784 9220 5840 9222
rect 6204 10906 6260 10908
rect 6284 10906 6340 10908
rect 6364 10906 6420 10908
rect 6444 10906 6500 10908
rect 6204 10854 6250 10906
rect 6250 10854 6260 10906
rect 6284 10854 6314 10906
rect 6314 10854 6326 10906
rect 6326 10854 6340 10906
rect 6364 10854 6378 10906
rect 6378 10854 6390 10906
rect 6390 10854 6420 10906
rect 6444 10854 6454 10906
rect 6454 10854 6500 10906
rect 6204 10852 6260 10854
rect 6284 10852 6340 10854
rect 6364 10852 6420 10854
rect 6444 10852 6500 10854
rect 6204 9818 6260 9820
rect 6284 9818 6340 9820
rect 6364 9818 6420 9820
rect 6444 9818 6500 9820
rect 6204 9766 6250 9818
rect 6250 9766 6260 9818
rect 6284 9766 6314 9818
rect 6314 9766 6326 9818
rect 6326 9766 6340 9818
rect 6364 9766 6378 9818
rect 6378 9766 6390 9818
rect 6390 9766 6420 9818
rect 6444 9766 6454 9818
rect 6454 9766 6500 9818
rect 6204 9764 6260 9766
rect 6284 9764 6340 9766
rect 6364 9764 6420 9766
rect 6444 9764 6500 9766
rect 9263 13082 9319 13084
rect 9343 13082 9399 13084
rect 9423 13082 9479 13084
rect 9503 13082 9559 13084
rect 9263 13030 9309 13082
rect 9309 13030 9319 13082
rect 9343 13030 9373 13082
rect 9373 13030 9385 13082
rect 9385 13030 9399 13082
rect 9423 13030 9437 13082
rect 9437 13030 9449 13082
rect 9449 13030 9479 13082
rect 9503 13030 9513 13082
rect 9513 13030 9559 13082
rect 9263 13028 9319 13030
rect 9343 13028 9399 13030
rect 9423 13028 9479 13030
rect 9503 13028 9559 13030
rect 8603 12538 8659 12540
rect 8683 12538 8739 12540
rect 8763 12538 8819 12540
rect 8843 12538 8899 12540
rect 8603 12486 8649 12538
rect 8649 12486 8659 12538
rect 8683 12486 8713 12538
rect 8713 12486 8725 12538
rect 8725 12486 8739 12538
rect 8763 12486 8777 12538
rect 8777 12486 8789 12538
rect 8789 12486 8819 12538
rect 8843 12486 8853 12538
rect 8853 12486 8899 12538
rect 8603 12484 8659 12486
rect 8683 12484 8739 12486
rect 8763 12484 8819 12486
rect 8843 12484 8899 12486
rect 8390 12164 8446 12200
rect 8390 12144 8392 12164
rect 8392 12144 8444 12164
rect 8444 12144 8446 12164
rect 8603 11450 8659 11452
rect 8683 11450 8739 11452
rect 8763 11450 8819 11452
rect 8843 11450 8899 11452
rect 8603 11398 8649 11450
rect 8649 11398 8659 11450
rect 8683 11398 8713 11450
rect 8713 11398 8725 11450
rect 8725 11398 8739 11450
rect 8763 11398 8777 11450
rect 8777 11398 8789 11450
rect 8789 11398 8819 11450
rect 8843 11398 8853 11450
rect 8853 11398 8899 11450
rect 8603 11396 8659 11398
rect 8683 11396 8739 11398
rect 8763 11396 8819 11398
rect 8843 11396 8899 11398
rect 9678 12044 9686 12064
rect 9686 12044 9734 12064
rect 9678 12008 9734 12044
rect 9263 11994 9319 11996
rect 9343 11994 9399 11996
rect 9423 11994 9479 11996
rect 9503 11994 9559 11996
rect 9263 11942 9309 11994
rect 9309 11942 9319 11994
rect 9343 11942 9373 11994
rect 9373 11942 9385 11994
rect 9385 11942 9399 11994
rect 9423 11942 9437 11994
rect 9437 11942 9449 11994
rect 9449 11942 9479 11994
rect 9503 11942 9513 11994
rect 9513 11942 9559 11994
rect 9263 11940 9319 11942
rect 9343 11940 9399 11942
rect 9423 11940 9479 11942
rect 9503 11940 9559 11942
rect 10138 12008 10194 12064
rect 11662 13626 11718 13628
rect 11742 13626 11798 13628
rect 11822 13626 11878 13628
rect 11902 13626 11958 13628
rect 11662 13574 11708 13626
rect 11708 13574 11718 13626
rect 11742 13574 11772 13626
rect 11772 13574 11784 13626
rect 11784 13574 11798 13626
rect 11822 13574 11836 13626
rect 11836 13574 11848 13626
rect 11848 13574 11878 13626
rect 11902 13574 11912 13626
rect 11912 13574 11958 13626
rect 11662 13572 11718 13574
rect 11742 13572 11798 13574
rect 11822 13572 11878 13574
rect 11902 13572 11958 13574
rect 11662 12538 11718 12540
rect 11742 12538 11798 12540
rect 11822 12538 11878 12540
rect 11902 12538 11958 12540
rect 11662 12486 11708 12538
rect 11708 12486 11718 12538
rect 11742 12486 11772 12538
rect 11772 12486 11784 12538
rect 11784 12486 11798 12538
rect 11822 12486 11836 12538
rect 11836 12486 11848 12538
rect 11848 12486 11878 12538
rect 11902 12486 11912 12538
rect 11912 12486 11958 12538
rect 11662 12484 11718 12486
rect 11742 12484 11798 12486
rect 11822 12484 11878 12486
rect 11902 12484 11958 12486
rect 12322 13082 12378 13084
rect 12402 13082 12458 13084
rect 12482 13082 12538 13084
rect 12562 13082 12618 13084
rect 12322 13030 12368 13082
rect 12368 13030 12378 13082
rect 12402 13030 12432 13082
rect 12432 13030 12444 13082
rect 12444 13030 12458 13082
rect 12482 13030 12496 13082
rect 12496 13030 12508 13082
rect 12508 13030 12538 13082
rect 12562 13030 12572 13082
rect 12572 13030 12618 13082
rect 12322 13028 12378 13030
rect 12402 13028 12458 13030
rect 12482 13028 12538 13030
rect 12562 13028 12618 13030
rect 9263 10906 9319 10908
rect 9343 10906 9399 10908
rect 9423 10906 9479 10908
rect 9503 10906 9559 10908
rect 9263 10854 9309 10906
rect 9309 10854 9319 10906
rect 9343 10854 9373 10906
rect 9373 10854 9385 10906
rect 9385 10854 9399 10906
rect 9423 10854 9437 10906
rect 9437 10854 9449 10906
rect 9449 10854 9479 10906
rect 9503 10854 9513 10906
rect 9513 10854 9559 10906
rect 9263 10852 9319 10854
rect 9343 10852 9399 10854
rect 9423 10852 9479 10854
rect 9503 10852 9559 10854
rect 6204 8730 6260 8732
rect 6284 8730 6340 8732
rect 6364 8730 6420 8732
rect 6444 8730 6500 8732
rect 6204 8678 6250 8730
rect 6250 8678 6260 8730
rect 6284 8678 6314 8730
rect 6314 8678 6326 8730
rect 6326 8678 6340 8730
rect 6364 8678 6378 8730
rect 6378 8678 6390 8730
rect 6390 8678 6420 8730
rect 6444 8678 6454 8730
rect 6454 8678 6500 8730
rect 6204 8676 6260 8678
rect 6284 8676 6340 8678
rect 6364 8676 6420 8678
rect 6444 8676 6500 8678
rect 5544 8186 5600 8188
rect 5624 8186 5680 8188
rect 5704 8186 5760 8188
rect 5784 8186 5840 8188
rect 5544 8134 5590 8186
rect 5590 8134 5600 8186
rect 5624 8134 5654 8186
rect 5654 8134 5666 8186
rect 5666 8134 5680 8186
rect 5704 8134 5718 8186
rect 5718 8134 5730 8186
rect 5730 8134 5760 8186
rect 5784 8134 5794 8186
rect 5794 8134 5840 8186
rect 5544 8132 5600 8134
rect 5624 8132 5680 8134
rect 5704 8132 5760 8134
rect 5784 8132 5840 8134
rect 6204 7642 6260 7644
rect 6284 7642 6340 7644
rect 6364 7642 6420 7644
rect 6444 7642 6500 7644
rect 6204 7590 6250 7642
rect 6250 7590 6260 7642
rect 6284 7590 6314 7642
rect 6314 7590 6326 7642
rect 6326 7590 6340 7642
rect 6364 7590 6378 7642
rect 6378 7590 6390 7642
rect 6390 7590 6420 7642
rect 6444 7590 6454 7642
rect 6454 7590 6500 7642
rect 6204 7588 6260 7590
rect 6284 7588 6340 7590
rect 6364 7588 6420 7590
rect 6444 7588 6500 7590
rect 5544 7098 5600 7100
rect 5624 7098 5680 7100
rect 5704 7098 5760 7100
rect 5784 7098 5840 7100
rect 5544 7046 5590 7098
rect 5590 7046 5600 7098
rect 5624 7046 5654 7098
rect 5654 7046 5666 7098
rect 5666 7046 5680 7098
rect 5704 7046 5718 7098
rect 5718 7046 5730 7098
rect 5730 7046 5760 7098
rect 5784 7046 5794 7098
rect 5794 7046 5840 7098
rect 5544 7044 5600 7046
rect 5624 7044 5680 7046
rect 5704 7044 5760 7046
rect 5784 7044 5840 7046
rect 6204 6554 6260 6556
rect 6284 6554 6340 6556
rect 6364 6554 6420 6556
rect 6444 6554 6500 6556
rect 6204 6502 6250 6554
rect 6250 6502 6260 6554
rect 6284 6502 6314 6554
rect 6314 6502 6326 6554
rect 6326 6502 6340 6554
rect 6364 6502 6378 6554
rect 6378 6502 6390 6554
rect 6390 6502 6420 6554
rect 6444 6502 6454 6554
rect 6454 6502 6500 6554
rect 6204 6500 6260 6502
rect 6284 6500 6340 6502
rect 6364 6500 6420 6502
rect 6444 6500 6500 6502
rect 5544 6010 5600 6012
rect 5624 6010 5680 6012
rect 5704 6010 5760 6012
rect 5784 6010 5840 6012
rect 5544 5958 5590 6010
rect 5590 5958 5600 6010
rect 5624 5958 5654 6010
rect 5654 5958 5666 6010
rect 5666 5958 5680 6010
rect 5704 5958 5718 6010
rect 5718 5958 5730 6010
rect 5730 5958 5760 6010
rect 5784 5958 5794 6010
rect 5794 5958 5840 6010
rect 5544 5956 5600 5958
rect 5624 5956 5680 5958
rect 5704 5956 5760 5958
rect 5784 5956 5840 5958
rect 6204 5466 6260 5468
rect 6284 5466 6340 5468
rect 6364 5466 6420 5468
rect 6444 5466 6500 5468
rect 6204 5414 6250 5466
rect 6250 5414 6260 5466
rect 6284 5414 6314 5466
rect 6314 5414 6326 5466
rect 6326 5414 6340 5466
rect 6364 5414 6378 5466
rect 6378 5414 6390 5466
rect 6390 5414 6420 5466
rect 6444 5414 6454 5466
rect 6454 5414 6500 5466
rect 6204 5412 6260 5414
rect 6284 5412 6340 5414
rect 6364 5412 6420 5414
rect 6444 5412 6500 5414
rect 5544 4922 5600 4924
rect 5624 4922 5680 4924
rect 5704 4922 5760 4924
rect 5784 4922 5840 4924
rect 5544 4870 5590 4922
rect 5590 4870 5600 4922
rect 5624 4870 5654 4922
rect 5654 4870 5666 4922
rect 5666 4870 5680 4922
rect 5704 4870 5718 4922
rect 5718 4870 5730 4922
rect 5730 4870 5760 4922
rect 5784 4870 5794 4922
rect 5794 4870 5840 4922
rect 5544 4868 5600 4870
rect 5624 4868 5680 4870
rect 5704 4868 5760 4870
rect 5784 4868 5840 4870
rect 6204 4378 6260 4380
rect 6284 4378 6340 4380
rect 6364 4378 6420 4380
rect 6444 4378 6500 4380
rect 6204 4326 6250 4378
rect 6250 4326 6260 4378
rect 6284 4326 6314 4378
rect 6314 4326 6326 4378
rect 6326 4326 6340 4378
rect 6364 4326 6378 4378
rect 6378 4326 6390 4378
rect 6390 4326 6420 4378
rect 6444 4326 6454 4378
rect 6454 4326 6500 4378
rect 6204 4324 6260 4326
rect 6284 4324 6340 4326
rect 6364 4324 6420 4326
rect 6444 4324 6500 4326
rect 8603 10362 8659 10364
rect 8683 10362 8739 10364
rect 8763 10362 8819 10364
rect 8843 10362 8899 10364
rect 8603 10310 8649 10362
rect 8649 10310 8659 10362
rect 8683 10310 8713 10362
rect 8713 10310 8725 10362
rect 8725 10310 8739 10362
rect 8763 10310 8777 10362
rect 8777 10310 8789 10362
rect 8789 10310 8819 10362
rect 8843 10310 8853 10362
rect 8853 10310 8899 10362
rect 8603 10308 8659 10310
rect 8683 10308 8739 10310
rect 8763 10308 8819 10310
rect 8843 10308 8899 10310
rect 9263 9818 9319 9820
rect 9343 9818 9399 9820
rect 9423 9818 9479 9820
rect 9503 9818 9559 9820
rect 9263 9766 9309 9818
rect 9309 9766 9319 9818
rect 9343 9766 9373 9818
rect 9373 9766 9385 9818
rect 9385 9766 9399 9818
rect 9423 9766 9437 9818
rect 9437 9766 9449 9818
rect 9449 9766 9479 9818
rect 9503 9766 9513 9818
rect 9513 9766 9559 9818
rect 9263 9764 9319 9766
rect 9343 9764 9399 9766
rect 9423 9764 9479 9766
rect 9503 9764 9559 9766
rect 11058 12144 11114 12200
rect 11662 11450 11718 11452
rect 11742 11450 11798 11452
rect 11822 11450 11878 11452
rect 11902 11450 11958 11452
rect 11662 11398 11708 11450
rect 11708 11398 11718 11450
rect 11742 11398 11772 11450
rect 11772 11398 11784 11450
rect 11784 11398 11798 11450
rect 11822 11398 11836 11450
rect 11836 11398 11848 11450
rect 11848 11398 11878 11450
rect 11902 11398 11912 11450
rect 11912 11398 11958 11450
rect 11662 11396 11718 11398
rect 11742 11396 11798 11398
rect 11822 11396 11878 11398
rect 11902 11396 11958 11398
rect 12322 11994 12378 11996
rect 12402 11994 12458 11996
rect 12482 11994 12538 11996
rect 12562 11994 12618 11996
rect 12322 11942 12368 11994
rect 12368 11942 12378 11994
rect 12402 11942 12432 11994
rect 12432 11942 12444 11994
rect 12444 11942 12458 11994
rect 12482 11942 12496 11994
rect 12496 11942 12508 11994
rect 12508 11942 12538 11994
rect 12562 11942 12572 11994
rect 12572 11942 12618 11994
rect 12322 11940 12378 11942
rect 12402 11940 12458 11942
rect 12482 11940 12538 11942
rect 12562 11940 12618 11942
rect 11662 10362 11718 10364
rect 11742 10362 11798 10364
rect 11822 10362 11878 10364
rect 11902 10362 11958 10364
rect 11662 10310 11708 10362
rect 11708 10310 11718 10362
rect 11742 10310 11772 10362
rect 11772 10310 11784 10362
rect 11784 10310 11798 10362
rect 11822 10310 11836 10362
rect 11836 10310 11848 10362
rect 11848 10310 11878 10362
rect 11902 10310 11912 10362
rect 11912 10310 11958 10362
rect 11662 10308 11718 10310
rect 11742 10308 11798 10310
rect 11822 10308 11878 10310
rect 11902 10308 11958 10310
rect 12322 10906 12378 10908
rect 12402 10906 12458 10908
rect 12482 10906 12538 10908
rect 12562 10906 12618 10908
rect 12322 10854 12368 10906
rect 12368 10854 12378 10906
rect 12402 10854 12432 10906
rect 12432 10854 12444 10906
rect 12444 10854 12458 10906
rect 12482 10854 12496 10906
rect 12496 10854 12508 10906
rect 12508 10854 12538 10906
rect 12562 10854 12572 10906
rect 12572 10854 12618 10906
rect 12322 10852 12378 10854
rect 12402 10852 12458 10854
rect 12482 10852 12538 10854
rect 12562 10852 12618 10854
rect 8603 9274 8659 9276
rect 8683 9274 8739 9276
rect 8763 9274 8819 9276
rect 8843 9274 8899 9276
rect 8603 9222 8649 9274
rect 8649 9222 8659 9274
rect 8683 9222 8713 9274
rect 8713 9222 8725 9274
rect 8725 9222 8739 9274
rect 8763 9222 8777 9274
rect 8777 9222 8789 9274
rect 8789 9222 8819 9274
rect 8843 9222 8853 9274
rect 8853 9222 8899 9274
rect 8603 9220 8659 9222
rect 8683 9220 8739 9222
rect 8763 9220 8819 9222
rect 8843 9220 8899 9222
rect 9263 8730 9319 8732
rect 9343 8730 9399 8732
rect 9423 8730 9479 8732
rect 9503 8730 9559 8732
rect 9263 8678 9309 8730
rect 9309 8678 9319 8730
rect 9343 8678 9373 8730
rect 9373 8678 9385 8730
rect 9385 8678 9399 8730
rect 9423 8678 9437 8730
rect 9437 8678 9449 8730
rect 9449 8678 9479 8730
rect 9503 8678 9513 8730
rect 9513 8678 9559 8730
rect 9263 8676 9319 8678
rect 9343 8676 9399 8678
rect 9423 8676 9479 8678
rect 9503 8676 9559 8678
rect 11662 9274 11718 9276
rect 11742 9274 11798 9276
rect 11822 9274 11878 9276
rect 11902 9274 11958 9276
rect 11662 9222 11708 9274
rect 11708 9222 11718 9274
rect 11742 9222 11772 9274
rect 11772 9222 11784 9274
rect 11784 9222 11798 9274
rect 11822 9222 11836 9274
rect 11836 9222 11848 9274
rect 11848 9222 11878 9274
rect 11902 9222 11912 9274
rect 11912 9222 11958 9274
rect 11662 9220 11718 9222
rect 11742 9220 11798 9222
rect 11822 9220 11878 9222
rect 11902 9220 11958 9222
rect 8603 8186 8659 8188
rect 8683 8186 8739 8188
rect 8763 8186 8819 8188
rect 8843 8186 8899 8188
rect 8603 8134 8649 8186
rect 8649 8134 8659 8186
rect 8683 8134 8713 8186
rect 8713 8134 8725 8186
rect 8725 8134 8739 8186
rect 8763 8134 8777 8186
rect 8777 8134 8789 8186
rect 8789 8134 8819 8186
rect 8843 8134 8853 8186
rect 8853 8134 8899 8186
rect 8603 8132 8659 8134
rect 8683 8132 8739 8134
rect 8763 8132 8819 8134
rect 8843 8132 8899 8134
rect 11662 8186 11718 8188
rect 11742 8186 11798 8188
rect 11822 8186 11878 8188
rect 11902 8186 11958 8188
rect 11662 8134 11708 8186
rect 11708 8134 11718 8186
rect 11742 8134 11772 8186
rect 11772 8134 11784 8186
rect 11784 8134 11798 8186
rect 11822 8134 11836 8186
rect 11836 8134 11848 8186
rect 11848 8134 11878 8186
rect 11902 8134 11912 8186
rect 11912 8134 11958 8186
rect 11662 8132 11718 8134
rect 11742 8132 11798 8134
rect 11822 8132 11878 8134
rect 11902 8132 11958 8134
rect 8603 7098 8659 7100
rect 8683 7098 8739 7100
rect 8763 7098 8819 7100
rect 8843 7098 8899 7100
rect 8603 7046 8649 7098
rect 8649 7046 8659 7098
rect 8683 7046 8713 7098
rect 8713 7046 8725 7098
rect 8725 7046 8739 7098
rect 8763 7046 8777 7098
rect 8777 7046 8789 7098
rect 8789 7046 8819 7098
rect 8843 7046 8853 7098
rect 8853 7046 8899 7098
rect 8603 7044 8659 7046
rect 8683 7044 8739 7046
rect 8763 7044 8819 7046
rect 8843 7044 8899 7046
rect 9263 7642 9319 7644
rect 9343 7642 9399 7644
rect 9423 7642 9479 7644
rect 9503 7642 9559 7644
rect 9263 7590 9309 7642
rect 9309 7590 9319 7642
rect 9343 7590 9373 7642
rect 9373 7590 9385 7642
rect 9385 7590 9399 7642
rect 9423 7590 9437 7642
rect 9437 7590 9449 7642
rect 9449 7590 9479 7642
rect 9503 7590 9513 7642
rect 9513 7590 9559 7642
rect 9263 7588 9319 7590
rect 9343 7588 9399 7590
rect 9423 7588 9479 7590
rect 9503 7588 9559 7590
rect 8603 6010 8659 6012
rect 8683 6010 8739 6012
rect 8763 6010 8819 6012
rect 8843 6010 8899 6012
rect 8603 5958 8649 6010
rect 8649 5958 8659 6010
rect 8683 5958 8713 6010
rect 8713 5958 8725 6010
rect 8725 5958 8739 6010
rect 8763 5958 8777 6010
rect 8777 5958 8789 6010
rect 8789 5958 8819 6010
rect 8843 5958 8853 6010
rect 8853 5958 8899 6010
rect 8603 5956 8659 5958
rect 8683 5956 8739 5958
rect 8763 5956 8819 5958
rect 8843 5956 8899 5958
rect 9263 6554 9319 6556
rect 9343 6554 9399 6556
rect 9423 6554 9479 6556
rect 9503 6554 9559 6556
rect 9263 6502 9309 6554
rect 9309 6502 9319 6554
rect 9343 6502 9373 6554
rect 9373 6502 9385 6554
rect 9385 6502 9399 6554
rect 9423 6502 9437 6554
rect 9437 6502 9449 6554
rect 9449 6502 9479 6554
rect 9503 6502 9513 6554
rect 9513 6502 9559 6554
rect 9263 6500 9319 6502
rect 9343 6500 9399 6502
rect 9423 6500 9479 6502
rect 9503 6500 9559 6502
rect 9263 5466 9319 5468
rect 9343 5466 9399 5468
rect 9423 5466 9479 5468
rect 9503 5466 9559 5468
rect 9263 5414 9309 5466
rect 9309 5414 9319 5466
rect 9343 5414 9373 5466
rect 9373 5414 9385 5466
rect 9385 5414 9399 5466
rect 9423 5414 9437 5466
rect 9437 5414 9449 5466
rect 9449 5414 9479 5466
rect 9503 5414 9513 5466
rect 9513 5414 9559 5466
rect 9263 5412 9319 5414
rect 9343 5412 9399 5414
rect 9423 5412 9479 5414
rect 9503 5412 9559 5414
rect 5446 4004 5502 4040
rect 5446 3984 5448 4004
rect 5448 3984 5500 4004
rect 5500 3984 5502 4004
rect 5544 3834 5600 3836
rect 5624 3834 5680 3836
rect 5704 3834 5760 3836
rect 5784 3834 5840 3836
rect 5544 3782 5590 3834
rect 5590 3782 5600 3834
rect 5624 3782 5654 3834
rect 5654 3782 5666 3834
rect 5666 3782 5680 3834
rect 5704 3782 5718 3834
rect 5718 3782 5730 3834
rect 5730 3782 5760 3834
rect 5784 3782 5794 3834
rect 5794 3782 5840 3834
rect 5544 3780 5600 3782
rect 5624 3780 5680 3782
rect 5704 3780 5760 3782
rect 5784 3780 5840 3782
rect 6458 3848 6514 3904
rect 6204 3290 6260 3292
rect 6284 3290 6340 3292
rect 6364 3290 6420 3292
rect 6444 3290 6500 3292
rect 6204 3238 6250 3290
rect 6250 3238 6260 3290
rect 6284 3238 6314 3290
rect 6314 3238 6326 3290
rect 6326 3238 6340 3290
rect 6364 3238 6378 3290
rect 6378 3238 6390 3290
rect 6390 3238 6420 3290
rect 6444 3238 6454 3290
rect 6454 3238 6500 3290
rect 6204 3236 6260 3238
rect 6284 3236 6340 3238
rect 6364 3236 6420 3238
rect 6444 3236 6500 3238
rect 7194 3476 7196 3496
rect 7196 3476 7248 3496
rect 7248 3476 7250 3496
rect 7194 3440 7250 3476
rect 5544 2746 5600 2748
rect 5624 2746 5680 2748
rect 5704 2746 5760 2748
rect 5784 2746 5840 2748
rect 5544 2694 5590 2746
rect 5590 2694 5600 2746
rect 5624 2694 5654 2746
rect 5654 2694 5666 2746
rect 5666 2694 5680 2746
rect 5704 2694 5718 2746
rect 5718 2694 5730 2746
rect 5730 2694 5760 2746
rect 5784 2694 5794 2746
rect 5794 2694 5840 2746
rect 5544 2692 5600 2694
rect 5624 2692 5680 2694
rect 5704 2692 5760 2694
rect 5784 2692 5840 2694
rect 8603 4922 8659 4924
rect 8683 4922 8739 4924
rect 8763 4922 8819 4924
rect 8843 4922 8899 4924
rect 8603 4870 8649 4922
rect 8649 4870 8659 4922
rect 8683 4870 8713 4922
rect 8713 4870 8725 4922
rect 8725 4870 8739 4922
rect 8763 4870 8777 4922
rect 8777 4870 8789 4922
rect 8789 4870 8819 4922
rect 8843 4870 8853 4922
rect 8853 4870 8899 4922
rect 8603 4868 8659 4870
rect 8683 4868 8739 4870
rect 8763 4868 8819 4870
rect 8843 4868 8899 4870
rect 9263 4378 9319 4380
rect 9343 4378 9399 4380
rect 9423 4378 9479 4380
rect 9503 4378 9559 4380
rect 9263 4326 9309 4378
rect 9309 4326 9319 4378
rect 9343 4326 9373 4378
rect 9373 4326 9385 4378
rect 9385 4326 9399 4378
rect 9423 4326 9437 4378
rect 9437 4326 9449 4378
rect 9449 4326 9479 4378
rect 9503 4326 9513 4378
rect 9513 4326 9559 4378
rect 9263 4324 9319 4326
rect 9343 4324 9399 4326
rect 9423 4324 9479 4326
rect 9503 4324 9559 4326
rect 11662 7098 11718 7100
rect 11742 7098 11798 7100
rect 11822 7098 11878 7100
rect 11902 7098 11958 7100
rect 11662 7046 11708 7098
rect 11708 7046 11718 7098
rect 11742 7046 11772 7098
rect 11772 7046 11784 7098
rect 11784 7046 11798 7098
rect 11822 7046 11836 7098
rect 11836 7046 11848 7098
rect 11848 7046 11878 7098
rect 11902 7046 11912 7098
rect 11912 7046 11958 7098
rect 11662 7044 11718 7046
rect 11742 7044 11798 7046
rect 11822 7044 11878 7046
rect 11902 7044 11958 7046
rect 12990 10104 13046 10160
rect 12322 9818 12378 9820
rect 12402 9818 12458 9820
rect 12482 9818 12538 9820
rect 12562 9818 12618 9820
rect 12322 9766 12368 9818
rect 12368 9766 12378 9818
rect 12402 9766 12432 9818
rect 12432 9766 12444 9818
rect 12444 9766 12458 9818
rect 12482 9766 12496 9818
rect 12496 9766 12508 9818
rect 12508 9766 12538 9818
rect 12562 9766 12572 9818
rect 12572 9766 12618 9818
rect 12322 9764 12378 9766
rect 12402 9764 12458 9766
rect 12482 9764 12538 9766
rect 12562 9764 12618 9766
rect 12322 8730 12378 8732
rect 12402 8730 12458 8732
rect 12482 8730 12538 8732
rect 12562 8730 12618 8732
rect 12322 8678 12368 8730
rect 12368 8678 12378 8730
rect 12402 8678 12432 8730
rect 12432 8678 12444 8730
rect 12444 8678 12458 8730
rect 12482 8678 12496 8730
rect 12496 8678 12508 8730
rect 12508 8678 12538 8730
rect 12562 8678 12572 8730
rect 12572 8678 12618 8730
rect 12322 8676 12378 8678
rect 12402 8676 12458 8678
rect 12482 8676 12538 8678
rect 12562 8676 12618 8678
rect 12322 7642 12378 7644
rect 12402 7642 12458 7644
rect 12482 7642 12538 7644
rect 12562 7642 12618 7644
rect 12322 7590 12368 7642
rect 12368 7590 12378 7642
rect 12402 7590 12432 7642
rect 12432 7590 12444 7642
rect 12444 7590 12458 7642
rect 12482 7590 12496 7642
rect 12496 7590 12508 7642
rect 12508 7590 12538 7642
rect 12562 7590 12572 7642
rect 12572 7590 12618 7642
rect 12322 7588 12378 7590
rect 12402 7588 12458 7590
rect 12482 7588 12538 7590
rect 12562 7588 12618 7590
rect 12322 6554 12378 6556
rect 12402 6554 12458 6556
rect 12482 6554 12538 6556
rect 12562 6554 12618 6556
rect 12322 6502 12368 6554
rect 12368 6502 12378 6554
rect 12402 6502 12432 6554
rect 12432 6502 12444 6554
rect 12444 6502 12458 6554
rect 12482 6502 12496 6554
rect 12496 6502 12508 6554
rect 12508 6502 12538 6554
rect 12562 6502 12572 6554
rect 12572 6502 12618 6554
rect 12322 6500 12378 6502
rect 12402 6500 12458 6502
rect 12482 6500 12538 6502
rect 12562 6500 12618 6502
rect 12990 6024 13046 6080
rect 11662 6010 11718 6012
rect 11742 6010 11798 6012
rect 11822 6010 11878 6012
rect 11902 6010 11958 6012
rect 11662 5958 11708 6010
rect 11708 5958 11718 6010
rect 11742 5958 11772 6010
rect 11772 5958 11784 6010
rect 11784 5958 11798 6010
rect 11822 5958 11836 6010
rect 11836 5958 11848 6010
rect 11848 5958 11878 6010
rect 11902 5958 11912 6010
rect 11912 5958 11958 6010
rect 11662 5956 11718 5958
rect 11742 5956 11798 5958
rect 11822 5956 11878 5958
rect 11902 5956 11958 5958
rect 12322 5466 12378 5468
rect 12402 5466 12458 5468
rect 12482 5466 12538 5468
rect 12562 5466 12618 5468
rect 12322 5414 12368 5466
rect 12368 5414 12378 5466
rect 12402 5414 12432 5466
rect 12432 5414 12444 5466
rect 12444 5414 12458 5466
rect 12482 5414 12496 5466
rect 12496 5414 12508 5466
rect 12508 5414 12538 5466
rect 12562 5414 12572 5466
rect 12572 5414 12618 5466
rect 12322 5412 12378 5414
rect 12402 5412 12458 5414
rect 12482 5412 12538 5414
rect 12562 5412 12618 5414
rect 8298 3848 8354 3904
rect 8603 3834 8659 3836
rect 8683 3834 8739 3836
rect 8763 3834 8819 3836
rect 8843 3834 8899 3836
rect 8603 3782 8649 3834
rect 8649 3782 8659 3834
rect 8683 3782 8713 3834
rect 8713 3782 8725 3834
rect 8725 3782 8739 3834
rect 8763 3782 8777 3834
rect 8777 3782 8789 3834
rect 8789 3782 8819 3834
rect 8843 3782 8853 3834
rect 8853 3782 8899 3834
rect 8603 3780 8659 3782
rect 8683 3780 8739 3782
rect 8763 3780 8819 3782
rect 8843 3780 8899 3782
rect 8298 3440 8354 3496
rect 9263 3290 9319 3292
rect 9343 3290 9399 3292
rect 9423 3290 9479 3292
rect 9503 3290 9559 3292
rect 9263 3238 9309 3290
rect 9309 3238 9319 3290
rect 9343 3238 9373 3290
rect 9373 3238 9385 3290
rect 9385 3238 9399 3290
rect 9423 3238 9437 3290
rect 9437 3238 9449 3290
rect 9449 3238 9479 3290
rect 9503 3238 9513 3290
rect 9513 3238 9559 3290
rect 9263 3236 9319 3238
rect 9343 3236 9399 3238
rect 9423 3236 9479 3238
rect 9503 3236 9559 3238
rect 11662 4922 11718 4924
rect 11742 4922 11798 4924
rect 11822 4922 11878 4924
rect 11902 4922 11958 4924
rect 11662 4870 11708 4922
rect 11708 4870 11718 4922
rect 11742 4870 11772 4922
rect 11772 4870 11784 4922
rect 11784 4870 11798 4922
rect 11822 4870 11836 4922
rect 11836 4870 11848 4922
rect 11848 4870 11878 4922
rect 11902 4870 11912 4922
rect 11912 4870 11958 4922
rect 11662 4868 11718 4870
rect 11742 4868 11798 4870
rect 11822 4868 11878 4870
rect 11902 4868 11958 4870
rect 12322 4378 12378 4380
rect 12402 4378 12458 4380
rect 12482 4378 12538 4380
rect 12562 4378 12618 4380
rect 12322 4326 12368 4378
rect 12368 4326 12378 4378
rect 12402 4326 12432 4378
rect 12432 4326 12444 4378
rect 12444 4326 12458 4378
rect 12482 4326 12496 4378
rect 12496 4326 12508 4378
rect 12508 4326 12538 4378
rect 12562 4326 12572 4378
rect 12572 4326 12618 4378
rect 12322 4324 12378 4326
rect 12402 4324 12458 4326
rect 12482 4324 12538 4326
rect 12562 4324 12618 4326
rect 11662 3834 11718 3836
rect 11742 3834 11798 3836
rect 11822 3834 11878 3836
rect 11902 3834 11958 3836
rect 11662 3782 11708 3834
rect 11708 3782 11718 3834
rect 11742 3782 11772 3834
rect 11772 3782 11784 3834
rect 11784 3782 11798 3834
rect 11822 3782 11836 3834
rect 11836 3782 11848 3834
rect 11848 3782 11878 3834
rect 11902 3782 11912 3834
rect 11912 3782 11958 3834
rect 11662 3780 11718 3782
rect 11742 3780 11798 3782
rect 11822 3780 11878 3782
rect 11902 3780 11958 3782
rect 8603 2746 8659 2748
rect 8683 2746 8739 2748
rect 8763 2746 8819 2748
rect 8843 2746 8899 2748
rect 8603 2694 8649 2746
rect 8649 2694 8659 2746
rect 8683 2694 8713 2746
rect 8713 2694 8725 2746
rect 8725 2694 8739 2746
rect 8763 2694 8777 2746
rect 8777 2694 8789 2746
rect 8789 2694 8819 2746
rect 8843 2694 8853 2746
rect 8853 2694 8899 2746
rect 8603 2692 8659 2694
rect 8683 2692 8739 2694
rect 8763 2692 8819 2694
rect 8843 2692 8899 2694
rect 12322 3290 12378 3292
rect 12402 3290 12458 3292
rect 12482 3290 12538 3292
rect 12562 3290 12618 3292
rect 12322 3238 12368 3290
rect 12368 3238 12378 3290
rect 12402 3238 12432 3290
rect 12432 3238 12444 3290
rect 12444 3238 12458 3290
rect 12482 3238 12496 3290
rect 12496 3238 12508 3290
rect 12508 3238 12538 3290
rect 12562 3238 12572 3290
rect 12572 3238 12618 3290
rect 12322 3236 12378 3238
rect 12402 3236 12458 3238
rect 12482 3236 12538 3238
rect 12562 3236 12618 3238
rect 11662 2746 11718 2748
rect 11742 2746 11798 2748
rect 11822 2746 11878 2748
rect 11902 2746 11958 2748
rect 11662 2694 11708 2746
rect 11708 2694 11718 2746
rect 11742 2694 11772 2746
rect 11772 2694 11784 2746
rect 11784 2694 11798 2746
rect 11822 2694 11836 2746
rect 11836 2694 11848 2746
rect 11848 2694 11878 2746
rect 11902 2694 11912 2746
rect 11912 2694 11958 2746
rect 11662 2692 11718 2694
rect 11742 2692 11798 2694
rect 11822 2692 11878 2694
rect 11902 2692 11958 2694
rect 3145 2202 3201 2204
rect 3225 2202 3281 2204
rect 3305 2202 3361 2204
rect 3385 2202 3441 2204
rect 3145 2150 3191 2202
rect 3191 2150 3201 2202
rect 3225 2150 3255 2202
rect 3255 2150 3267 2202
rect 3267 2150 3281 2202
rect 3305 2150 3319 2202
rect 3319 2150 3331 2202
rect 3331 2150 3361 2202
rect 3385 2150 3395 2202
rect 3395 2150 3441 2202
rect 3145 2148 3201 2150
rect 3225 2148 3281 2150
rect 3305 2148 3361 2150
rect 3385 2148 3441 2150
rect 6204 2202 6260 2204
rect 6284 2202 6340 2204
rect 6364 2202 6420 2204
rect 6444 2202 6500 2204
rect 6204 2150 6250 2202
rect 6250 2150 6260 2202
rect 6284 2150 6314 2202
rect 6314 2150 6326 2202
rect 6326 2150 6340 2202
rect 6364 2150 6378 2202
rect 6378 2150 6390 2202
rect 6390 2150 6420 2202
rect 6444 2150 6454 2202
rect 6454 2150 6500 2202
rect 6204 2148 6260 2150
rect 6284 2148 6340 2150
rect 6364 2148 6420 2150
rect 6444 2148 6500 2150
rect 9263 2202 9319 2204
rect 9343 2202 9399 2204
rect 9423 2202 9479 2204
rect 9503 2202 9559 2204
rect 9263 2150 9309 2202
rect 9309 2150 9319 2202
rect 9343 2150 9373 2202
rect 9373 2150 9385 2202
rect 9385 2150 9399 2202
rect 9423 2150 9437 2202
rect 9437 2150 9449 2202
rect 9449 2150 9479 2202
rect 9503 2150 9513 2202
rect 9513 2150 9559 2202
rect 9263 2148 9319 2150
rect 9343 2148 9399 2150
rect 9423 2148 9479 2150
rect 9503 2148 9559 2150
rect 12322 2202 12378 2204
rect 12402 2202 12458 2204
rect 12482 2202 12538 2204
rect 12562 2202 12618 2204
rect 12322 2150 12368 2202
rect 12368 2150 12378 2202
rect 12402 2150 12432 2202
rect 12432 2150 12444 2202
rect 12444 2150 12458 2202
rect 12482 2150 12496 2202
rect 12496 2150 12508 2202
rect 12508 2150 12538 2202
rect 12562 2150 12572 2202
rect 12572 2150 12618 2202
rect 12322 2148 12378 2150
rect 12402 2148 12458 2150
rect 12482 2148 12538 2150
rect 12562 2148 12618 2150
rect 13266 1944 13322 2000
<< metal3 >>
rect 13261 14242 13327 14245
rect 13657 14242 14457 14272
rect 13261 14240 14457 14242
rect 13261 14184 13266 14240
rect 13322 14184 14457 14240
rect 13261 14182 14457 14184
rect 13261 14179 13327 14182
rect 3135 14176 3451 14177
rect 3135 14112 3141 14176
rect 3205 14112 3221 14176
rect 3285 14112 3301 14176
rect 3365 14112 3381 14176
rect 3445 14112 3451 14176
rect 3135 14111 3451 14112
rect 6194 14176 6510 14177
rect 6194 14112 6200 14176
rect 6264 14112 6280 14176
rect 6344 14112 6360 14176
rect 6424 14112 6440 14176
rect 6504 14112 6510 14176
rect 6194 14111 6510 14112
rect 9253 14176 9569 14177
rect 9253 14112 9259 14176
rect 9323 14112 9339 14176
rect 9403 14112 9419 14176
rect 9483 14112 9499 14176
rect 9563 14112 9569 14176
rect 9253 14111 9569 14112
rect 12312 14176 12628 14177
rect 12312 14112 12318 14176
rect 12382 14112 12398 14176
rect 12462 14112 12478 14176
rect 12542 14112 12558 14176
rect 12622 14112 12628 14176
rect 13657 14152 14457 14182
rect 12312 14111 12628 14112
rect 2475 13632 2791 13633
rect 2475 13568 2481 13632
rect 2545 13568 2561 13632
rect 2625 13568 2641 13632
rect 2705 13568 2721 13632
rect 2785 13568 2791 13632
rect 2475 13567 2791 13568
rect 5534 13632 5850 13633
rect 5534 13568 5540 13632
rect 5604 13568 5620 13632
rect 5684 13568 5700 13632
rect 5764 13568 5780 13632
rect 5844 13568 5850 13632
rect 5534 13567 5850 13568
rect 8593 13632 8909 13633
rect 8593 13568 8599 13632
rect 8663 13568 8679 13632
rect 8743 13568 8759 13632
rect 8823 13568 8839 13632
rect 8903 13568 8909 13632
rect 8593 13567 8909 13568
rect 11652 13632 11968 13633
rect 11652 13568 11658 13632
rect 11722 13568 11738 13632
rect 11802 13568 11818 13632
rect 11882 13568 11898 13632
rect 11962 13568 11968 13632
rect 11652 13567 11968 13568
rect 3135 13088 3451 13089
rect 3135 13024 3141 13088
rect 3205 13024 3221 13088
rect 3285 13024 3301 13088
rect 3365 13024 3381 13088
rect 3445 13024 3451 13088
rect 3135 13023 3451 13024
rect 6194 13088 6510 13089
rect 6194 13024 6200 13088
rect 6264 13024 6280 13088
rect 6344 13024 6360 13088
rect 6424 13024 6440 13088
rect 6504 13024 6510 13088
rect 6194 13023 6510 13024
rect 9253 13088 9569 13089
rect 9253 13024 9259 13088
rect 9323 13024 9339 13088
rect 9403 13024 9419 13088
rect 9483 13024 9499 13088
rect 9563 13024 9569 13088
rect 9253 13023 9569 13024
rect 12312 13088 12628 13089
rect 12312 13024 12318 13088
rect 12382 13024 12398 13088
rect 12462 13024 12478 13088
rect 12542 13024 12558 13088
rect 12622 13024 12628 13088
rect 12312 13023 12628 13024
rect 2475 12544 2791 12545
rect 2475 12480 2481 12544
rect 2545 12480 2561 12544
rect 2625 12480 2641 12544
rect 2705 12480 2721 12544
rect 2785 12480 2791 12544
rect 2475 12479 2791 12480
rect 5534 12544 5850 12545
rect 5534 12480 5540 12544
rect 5604 12480 5620 12544
rect 5684 12480 5700 12544
rect 5764 12480 5780 12544
rect 5844 12480 5850 12544
rect 5534 12479 5850 12480
rect 8593 12544 8909 12545
rect 8593 12480 8599 12544
rect 8663 12480 8679 12544
rect 8743 12480 8759 12544
rect 8823 12480 8839 12544
rect 8903 12480 8909 12544
rect 8593 12479 8909 12480
rect 11652 12544 11968 12545
rect 11652 12480 11658 12544
rect 11722 12480 11738 12544
rect 11802 12480 11818 12544
rect 11882 12480 11898 12544
rect 11962 12480 11968 12544
rect 11652 12479 11968 12480
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 8385 12202 8451 12205
rect 11053 12202 11119 12205
rect 8385 12200 11119 12202
rect 8385 12144 8390 12200
rect 8446 12144 11058 12200
rect 11114 12144 11119 12200
rect 8385 12142 11119 12144
rect 8385 12139 8451 12142
rect 11053 12139 11119 12142
rect 9673 12066 9739 12069
rect 10133 12066 10199 12069
rect 9673 12064 10199 12066
rect 9673 12008 9678 12064
rect 9734 12008 10138 12064
rect 10194 12008 10199 12064
rect 9673 12006 10199 12008
rect 9673 12003 9739 12006
rect 10133 12003 10199 12006
rect 3135 12000 3451 12001
rect 3135 11936 3141 12000
rect 3205 11936 3221 12000
rect 3285 11936 3301 12000
rect 3365 11936 3381 12000
rect 3445 11936 3451 12000
rect 3135 11935 3451 11936
rect 6194 12000 6510 12001
rect 6194 11936 6200 12000
rect 6264 11936 6280 12000
rect 6344 11936 6360 12000
rect 6424 11936 6440 12000
rect 6504 11936 6510 12000
rect 6194 11935 6510 11936
rect 9253 12000 9569 12001
rect 9253 11936 9259 12000
rect 9323 11936 9339 12000
rect 9403 11936 9419 12000
rect 9483 11936 9499 12000
rect 9563 11936 9569 12000
rect 9253 11935 9569 11936
rect 12312 12000 12628 12001
rect 12312 11936 12318 12000
rect 12382 11936 12398 12000
rect 12462 11936 12478 12000
rect 12542 11936 12558 12000
rect 12622 11936 12628 12000
rect 12312 11935 12628 11936
rect 2475 11456 2791 11457
rect 2475 11392 2481 11456
rect 2545 11392 2561 11456
rect 2625 11392 2641 11456
rect 2705 11392 2721 11456
rect 2785 11392 2791 11456
rect 2475 11391 2791 11392
rect 5534 11456 5850 11457
rect 5534 11392 5540 11456
rect 5604 11392 5620 11456
rect 5684 11392 5700 11456
rect 5764 11392 5780 11456
rect 5844 11392 5850 11456
rect 5534 11391 5850 11392
rect 8593 11456 8909 11457
rect 8593 11392 8599 11456
rect 8663 11392 8679 11456
rect 8743 11392 8759 11456
rect 8823 11392 8839 11456
rect 8903 11392 8909 11456
rect 8593 11391 8909 11392
rect 11652 11456 11968 11457
rect 11652 11392 11658 11456
rect 11722 11392 11738 11456
rect 11802 11392 11818 11456
rect 11882 11392 11898 11456
rect 11962 11392 11968 11456
rect 11652 11391 11968 11392
rect 3135 10912 3451 10913
rect 3135 10848 3141 10912
rect 3205 10848 3221 10912
rect 3285 10848 3301 10912
rect 3365 10848 3381 10912
rect 3445 10848 3451 10912
rect 3135 10847 3451 10848
rect 6194 10912 6510 10913
rect 6194 10848 6200 10912
rect 6264 10848 6280 10912
rect 6344 10848 6360 10912
rect 6424 10848 6440 10912
rect 6504 10848 6510 10912
rect 6194 10847 6510 10848
rect 9253 10912 9569 10913
rect 9253 10848 9259 10912
rect 9323 10848 9339 10912
rect 9403 10848 9419 10912
rect 9483 10848 9499 10912
rect 9563 10848 9569 10912
rect 9253 10847 9569 10848
rect 12312 10912 12628 10913
rect 12312 10848 12318 10912
rect 12382 10848 12398 10912
rect 12462 10848 12478 10912
rect 12542 10848 12558 10912
rect 12622 10848 12628 10912
rect 12312 10847 12628 10848
rect 2475 10368 2791 10369
rect 2475 10304 2481 10368
rect 2545 10304 2561 10368
rect 2625 10304 2641 10368
rect 2705 10304 2721 10368
rect 2785 10304 2791 10368
rect 2475 10303 2791 10304
rect 5534 10368 5850 10369
rect 5534 10304 5540 10368
rect 5604 10304 5620 10368
rect 5684 10304 5700 10368
rect 5764 10304 5780 10368
rect 5844 10304 5850 10368
rect 5534 10303 5850 10304
rect 8593 10368 8909 10369
rect 8593 10304 8599 10368
rect 8663 10304 8679 10368
rect 8743 10304 8759 10368
rect 8823 10304 8839 10368
rect 8903 10304 8909 10368
rect 8593 10303 8909 10304
rect 11652 10368 11968 10369
rect 11652 10304 11658 10368
rect 11722 10304 11738 10368
rect 11802 10304 11818 10368
rect 11882 10304 11898 10368
rect 11962 10304 11968 10368
rect 11652 10303 11968 10304
rect 12985 10162 13051 10165
rect 13657 10162 14457 10192
rect 12985 10160 14457 10162
rect 12985 10104 12990 10160
rect 13046 10104 14457 10160
rect 12985 10102 14457 10104
rect 12985 10099 13051 10102
rect 13657 10072 14457 10102
rect 3135 9824 3451 9825
rect 3135 9760 3141 9824
rect 3205 9760 3221 9824
rect 3285 9760 3301 9824
rect 3365 9760 3381 9824
rect 3445 9760 3451 9824
rect 3135 9759 3451 9760
rect 6194 9824 6510 9825
rect 6194 9760 6200 9824
rect 6264 9760 6280 9824
rect 6344 9760 6360 9824
rect 6424 9760 6440 9824
rect 6504 9760 6510 9824
rect 6194 9759 6510 9760
rect 9253 9824 9569 9825
rect 9253 9760 9259 9824
rect 9323 9760 9339 9824
rect 9403 9760 9419 9824
rect 9483 9760 9499 9824
rect 9563 9760 9569 9824
rect 9253 9759 9569 9760
rect 12312 9824 12628 9825
rect 12312 9760 12318 9824
rect 12382 9760 12398 9824
rect 12462 9760 12478 9824
rect 12542 9760 12558 9824
rect 12622 9760 12628 9824
rect 12312 9759 12628 9760
rect 2475 9280 2791 9281
rect 2475 9216 2481 9280
rect 2545 9216 2561 9280
rect 2625 9216 2641 9280
rect 2705 9216 2721 9280
rect 2785 9216 2791 9280
rect 2475 9215 2791 9216
rect 5534 9280 5850 9281
rect 5534 9216 5540 9280
rect 5604 9216 5620 9280
rect 5684 9216 5700 9280
rect 5764 9216 5780 9280
rect 5844 9216 5850 9280
rect 5534 9215 5850 9216
rect 8593 9280 8909 9281
rect 8593 9216 8599 9280
rect 8663 9216 8679 9280
rect 8743 9216 8759 9280
rect 8823 9216 8839 9280
rect 8903 9216 8909 9280
rect 8593 9215 8909 9216
rect 11652 9280 11968 9281
rect 11652 9216 11658 9280
rect 11722 9216 11738 9280
rect 11802 9216 11818 9280
rect 11882 9216 11898 9280
rect 11962 9216 11968 9280
rect 11652 9215 11968 9216
rect 3135 8736 3451 8737
rect 3135 8672 3141 8736
rect 3205 8672 3221 8736
rect 3285 8672 3301 8736
rect 3365 8672 3381 8736
rect 3445 8672 3451 8736
rect 3135 8671 3451 8672
rect 6194 8736 6510 8737
rect 6194 8672 6200 8736
rect 6264 8672 6280 8736
rect 6344 8672 6360 8736
rect 6424 8672 6440 8736
rect 6504 8672 6510 8736
rect 6194 8671 6510 8672
rect 9253 8736 9569 8737
rect 9253 8672 9259 8736
rect 9323 8672 9339 8736
rect 9403 8672 9419 8736
rect 9483 8672 9499 8736
rect 9563 8672 9569 8736
rect 9253 8671 9569 8672
rect 12312 8736 12628 8737
rect 12312 8672 12318 8736
rect 12382 8672 12398 8736
rect 12462 8672 12478 8736
rect 12542 8672 12558 8736
rect 12622 8672 12628 8736
rect 12312 8671 12628 8672
rect 2475 8192 2791 8193
rect 2475 8128 2481 8192
rect 2545 8128 2561 8192
rect 2625 8128 2641 8192
rect 2705 8128 2721 8192
rect 2785 8128 2791 8192
rect 2475 8127 2791 8128
rect 5534 8192 5850 8193
rect 5534 8128 5540 8192
rect 5604 8128 5620 8192
rect 5684 8128 5700 8192
rect 5764 8128 5780 8192
rect 5844 8128 5850 8192
rect 5534 8127 5850 8128
rect 8593 8192 8909 8193
rect 8593 8128 8599 8192
rect 8663 8128 8679 8192
rect 8743 8128 8759 8192
rect 8823 8128 8839 8192
rect 8903 8128 8909 8192
rect 8593 8127 8909 8128
rect 11652 8192 11968 8193
rect 11652 8128 11658 8192
rect 11722 8128 11738 8192
rect 11802 8128 11818 8192
rect 11882 8128 11898 8192
rect 11962 8128 11968 8192
rect 11652 8127 11968 8128
rect 3135 7648 3451 7649
rect 3135 7584 3141 7648
rect 3205 7584 3221 7648
rect 3285 7584 3301 7648
rect 3365 7584 3381 7648
rect 3445 7584 3451 7648
rect 3135 7583 3451 7584
rect 6194 7648 6510 7649
rect 6194 7584 6200 7648
rect 6264 7584 6280 7648
rect 6344 7584 6360 7648
rect 6424 7584 6440 7648
rect 6504 7584 6510 7648
rect 6194 7583 6510 7584
rect 9253 7648 9569 7649
rect 9253 7584 9259 7648
rect 9323 7584 9339 7648
rect 9403 7584 9419 7648
rect 9483 7584 9499 7648
rect 9563 7584 9569 7648
rect 9253 7583 9569 7584
rect 12312 7648 12628 7649
rect 12312 7584 12318 7648
rect 12382 7584 12398 7648
rect 12462 7584 12478 7648
rect 12542 7584 12558 7648
rect 12622 7584 12628 7648
rect 12312 7583 12628 7584
rect 2475 7104 2791 7105
rect 2475 7040 2481 7104
rect 2545 7040 2561 7104
rect 2625 7040 2641 7104
rect 2705 7040 2721 7104
rect 2785 7040 2791 7104
rect 2475 7039 2791 7040
rect 5534 7104 5850 7105
rect 5534 7040 5540 7104
rect 5604 7040 5620 7104
rect 5684 7040 5700 7104
rect 5764 7040 5780 7104
rect 5844 7040 5850 7104
rect 5534 7039 5850 7040
rect 8593 7104 8909 7105
rect 8593 7040 8599 7104
rect 8663 7040 8679 7104
rect 8743 7040 8759 7104
rect 8823 7040 8839 7104
rect 8903 7040 8909 7104
rect 8593 7039 8909 7040
rect 11652 7104 11968 7105
rect 11652 7040 11658 7104
rect 11722 7040 11738 7104
rect 11802 7040 11818 7104
rect 11882 7040 11898 7104
rect 11962 7040 11968 7104
rect 11652 7039 11968 7040
rect 3135 6560 3451 6561
rect 3135 6496 3141 6560
rect 3205 6496 3221 6560
rect 3285 6496 3301 6560
rect 3365 6496 3381 6560
rect 3445 6496 3451 6560
rect 3135 6495 3451 6496
rect 6194 6560 6510 6561
rect 6194 6496 6200 6560
rect 6264 6496 6280 6560
rect 6344 6496 6360 6560
rect 6424 6496 6440 6560
rect 6504 6496 6510 6560
rect 6194 6495 6510 6496
rect 9253 6560 9569 6561
rect 9253 6496 9259 6560
rect 9323 6496 9339 6560
rect 9403 6496 9419 6560
rect 9483 6496 9499 6560
rect 9563 6496 9569 6560
rect 9253 6495 9569 6496
rect 12312 6560 12628 6561
rect 12312 6496 12318 6560
rect 12382 6496 12398 6560
rect 12462 6496 12478 6560
rect 12542 6496 12558 6560
rect 12622 6496 12628 6560
rect 12312 6495 12628 6496
rect 12985 6082 13051 6085
rect 13657 6082 14457 6112
rect 12985 6080 14457 6082
rect 12985 6024 12990 6080
rect 13046 6024 14457 6080
rect 12985 6022 14457 6024
rect 12985 6019 13051 6022
rect 2475 6016 2791 6017
rect 2475 5952 2481 6016
rect 2545 5952 2561 6016
rect 2625 5952 2641 6016
rect 2705 5952 2721 6016
rect 2785 5952 2791 6016
rect 2475 5951 2791 5952
rect 5534 6016 5850 6017
rect 5534 5952 5540 6016
rect 5604 5952 5620 6016
rect 5684 5952 5700 6016
rect 5764 5952 5780 6016
rect 5844 5952 5850 6016
rect 5534 5951 5850 5952
rect 8593 6016 8909 6017
rect 8593 5952 8599 6016
rect 8663 5952 8679 6016
rect 8743 5952 8759 6016
rect 8823 5952 8839 6016
rect 8903 5952 8909 6016
rect 8593 5951 8909 5952
rect 11652 6016 11968 6017
rect 11652 5952 11658 6016
rect 11722 5952 11738 6016
rect 11802 5952 11818 6016
rect 11882 5952 11898 6016
rect 11962 5952 11968 6016
rect 13657 5992 14457 6022
rect 11652 5951 11968 5952
rect 3135 5472 3451 5473
rect 3135 5408 3141 5472
rect 3205 5408 3221 5472
rect 3285 5408 3301 5472
rect 3365 5408 3381 5472
rect 3445 5408 3451 5472
rect 3135 5407 3451 5408
rect 6194 5472 6510 5473
rect 6194 5408 6200 5472
rect 6264 5408 6280 5472
rect 6344 5408 6360 5472
rect 6424 5408 6440 5472
rect 6504 5408 6510 5472
rect 6194 5407 6510 5408
rect 9253 5472 9569 5473
rect 9253 5408 9259 5472
rect 9323 5408 9339 5472
rect 9403 5408 9419 5472
rect 9483 5408 9499 5472
rect 9563 5408 9569 5472
rect 9253 5407 9569 5408
rect 12312 5472 12628 5473
rect 12312 5408 12318 5472
rect 12382 5408 12398 5472
rect 12462 5408 12478 5472
rect 12542 5408 12558 5472
rect 12622 5408 12628 5472
rect 12312 5407 12628 5408
rect 2475 4928 2791 4929
rect 2475 4864 2481 4928
rect 2545 4864 2561 4928
rect 2625 4864 2641 4928
rect 2705 4864 2721 4928
rect 2785 4864 2791 4928
rect 2475 4863 2791 4864
rect 5534 4928 5850 4929
rect 5534 4864 5540 4928
rect 5604 4864 5620 4928
rect 5684 4864 5700 4928
rect 5764 4864 5780 4928
rect 5844 4864 5850 4928
rect 5534 4863 5850 4864
rect 8593 4928 8909 4929
rect 8593 4864 8599 4928
rect 8663 4864 8679 4928
rect 8743 4864 8759 4928
rect 8823 4864 8839 4928
rect 8903 4864 8909 4928
rect 8593 4863 8909 4864
rect 11652 4928 11968 4929
rect 11652 4864 11658 4928
rect 11722 4864 11738 4928
rect 11802 4864 11818 4928
rect 11882 4864 11898 4928
rect 11962 4864 11968 4928
rect 11652 4863 11968 4864
rect 3135 4384 3451 4385
rect 3135 4320 3141 4384
rect 3205 4320 3221 4384
rect 3285 4320 3301 4384
rect 3365 4320 3381 4384
rect 3445 4320 3451 4384
rect 3135 4319 3451 4320
rect 6194 4384 6510 4385
rect 6194 4320 6200 4384
rect 6264 4320 6280 4384
rect 6344 4320 6360 4384
rect 6424 4320 6440 4384
rect 6504 4320 6510 4384
rect 6194 4319 6510 4320
rect 9253 4384 9569 4385
rect 9253 4320 9259 4384
rect 9323 4320 9339 4384
rect 9403 4320 9419 4384
rect 9483 4320 9499 4384
rect 9563 4320 9569 4384
rect 9253 4319 9569 4320
rect 12312 4384 12628 4385
rect 12312 4320 12318 4384
rect 12382 4320 12398 4384
rect 12462 4320 12478 4384
rect 12542 4320 12558 4384
rect 12622 4320 12628 4384
rect 12312 4319 12628 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 2681 4042 2747 4045
rect 5441 4042 5507 4045
rect 2681 4040 5507 4042
rect 2681 3984 2686 4040
rect 2742 3984 5446 4040
rect 5502 3984 5507 4040
rect 2681 3982 5507 3984
rect 2681 3979 2747 3982
rect 5441 3979 5507 3982
rect 6453 3906 6519 3909
rect 8293 3906 8359 3909
rect 6453 3904 8359 3906
rect 6453 3848 6458 3904
rect 6514 3848 8298 3904
rect 8354 3848 8359 3904
rect 6453 3846 8359 3848
rect 6453 3843 6519 3846
rect 8293 3843 8359 3846
rect 2475 3840 2791 3841
rect 2475 3776 2481 3840
rect 2545 3776 2561 3840
rect 2625 3776 2641 3840
rect 2705 3776 2721 3840
rect 2785 3776 2791 3840
rect 2475 3775 2791 3776
rect 5534 3840 5850 3841
rect 5534 3776 5540 3840
rect 5604 3776 5620 3840
rect 5684 3776 5700 3840
rect 5764 3776 5780 3840
rect 5844 3776 5850 3840
rect 5534 3775 5850 3776
rect 8593 3840 8909 3841
rect 8593 3776 8599 3840
rect 8663 3776 8679 3840
rect 8743 3776 8759 3840
rect 8823 3776 8839 3840
rect 8903 3776 8909 3840
rect 8593 3775 8909 3776
rect 11652 3840 11968 3841
rect 11652 3776 11658 3840
rect 11722 3776 11738 3840
rect 11802 3776 11818 3840
rect 11882 3776 11898 3840
rect 11962 3776 11968 3840
rect 11652 3775 11968 3776
rect 7189 3498 7255 3501
rect 8293 3498 8359 3501
rect 7189 3496 8359 3498
rect 7189 3440 7194 3496
rect 7250 3440 8298 3496
rect 8354 3440 8359 3496
rect 7189 3438 8359 3440
rect 7189 3435 7255 3438
rect 8293 3435 8359 3438
rect 3135 3296 3451 3297
rect 3135 3232 3141 3296
rect 3205 3232 3221 3296
rect 3285 3232 3301 3296
rect 3365 3232 3381 3296
rect 3445 3232 3451 3296
rect 3135 3231 3451 3232
rect 6194 3296 6510 3297
rect 6194 3232 6200 3296
rect 6264 3232 6280 3296
rect 6344 3232 6360 3296
rect 6424 3232 6440 3296
rect 6504 3232 6510 3296
rect 6194 3231 6510 3232
rect 9253 3296 9569 3297
rect 9253 3232 9259 3296
rect 9323 3232 9339 3296
rect 9403 3232 9419 3296
rect 9483 3232 9499 3296
rect 9563 3232 9569 3296
rect 9253 3231 9569 3232
rect 12312 3296 12628 3297
rect 12312 3232 12318 3296
rect 12382 3232 12398 3296
rect 12462 3232 12478 3296
rect 12542 3232 12558 3296
rect 12622 3232 12628 3296
rect 12312 3231 12628 3232
rect 2475 2752 2791 2753
rect 2475 2688 2481 2752
rect 2545 2688 2561 2752
rect 2625 2688 2641 2752
rect 2705 2688 2721 2752
rect 2785 2688 2791 2752
rect 2475 2687 2791 2688
rect 5534 2752 5850 2753
rect 5534 2688 5540 2752
rect 5604 2688 5620 2752
rect 5684 2688 5700 2752
rect 5764 2688 5780 2752
rect 5844 2688 5850 2752
rect 5534 2687 5850 2688
rect 8593 2752 8909 2753
rect 8593 2688 8599 2752
rect 8663 2688 8679 2752
rect 8743 2688 8759 2752
rect 8823 2688 8839 2752
rect 8903 2688 8909 2752
rect 8593 2687 8909 2688
rect 11652 2752 11968 2753
rect 11652 2688 11658 2752
rect 11722 2688 11738 2752
rect 11802 2688 11818 2752
rect 11882 2688 11898 2752
rect 11962 2688 11968 2752
rect 11652 2687 11968 2688
rect 3135 2208 3451 2209
rect 3135 2144 3141 2208
rect 3205 2144 3221 2208
rect 3285 2144 3301 2208
rect 3365 2144 3381 2208
rect 3445 2144 3451 2208
rect 3135 2143 3451 2144
rect 6194 2208 6510 2209
rect 6194 2144 6200 2208
rect 6264 2144 6280 2208
rect 6344 2144 6360 2208
rect 6424 2144 6440 2208
rect 6504 2144 6510 2208
rect 6194 2143 6510 2144
rect 9253 2208 9569 2209
rect 9253 2144 9259 2208
rect 9323 2144 9339 2208
rect 9403 2144 9419 2208
rect 9483 2144 9499 2208
rect 9563 2144 9569 2208
rect 9253 2143 9569 2144
rect 12312 2208 12628 2209
rect 12312 2144 12318 2208
rect 12382 2144 12398 2208
rect 12462 2144 12478 2208
rect 12542 2144 12558 2208
rect 12622 2144 12628 2208
rect 12312 2143 12628 2144
rect 13261 2002 13327 2005
rect 13657 2002 14457 2032
rect 13261 2000 14457 2002
rect 13261 1944 13266 2000
rect 13322 1944 14457 2000
rect 13261 1942 14457 1944
rect 13261 1939 13327 1942
rect 13657 1912 14457 1942
<< via3 >>
rect 3141 14172 3205 14176
rect 3141 14116 3145 14172
rect 3145 14116 3201 14172
rect 3201 14116 3205 14172
rect 3141 14112 3205 14116
rect 3221 14172 3285 14176
rect 3221 14116 3225 14172
rect 3225 14116 3281 14172
rect 3281 14116 3285 14172
rect 3221 14112 3285 14116
rect 3301 14172 3365 14176
rect 3301 14116 3305 14172
rect 3305 14116 3361 14172
rect 3361 14116 3365 14172
rect 3301 14112 3365 14116
rect 3381 14172 3445 14176
rect 3381 14116 3385 14172
rect 3385 14116 3441 14172
rect 3441 14116 3445 14172
rect 3381 14112 3445 14116
rect 6200 14172 6264 14176
rect 6200 14116 6204 14172
rect 6204 14116 6260 14172
rect 6260 14116 6264 14172
rect 6200 14112 6264 14116
rect 6280 14172 6344 14176
rect 6280 14116 6284 14172
rect 6284 14116 6340 14172
rect 6340 14116 6344 14172
rect 6280 14112 6344 14116
rect 6360 14172 6424 14176
rect 6360 14116 6364 14172
rect 6364 14116 6420 14172
rect 6420 14116 6424 14172
rect 6360 14112 6424 14116
rect 6440 14172 6504 14176
rect 6440 14116 6444 14172
rect 6444 14116 6500 14172
rect 6500 14116 6504 14172
rect 6440 14112 6504 14116
rect 9259 14172 9323 14176
rect 9259 14116 9263 14172
rect 9263 14116 9319 14172
rect 9319 14116 9323 14172
rect 9259 14112 9323 14116
rect 9339 14172 9403 14176
rect 9339 14116 9343 14172
rect 9343 14116 9399 14172
rect 9399 14116 9403 14172
rect 9339 14112 9403 14116
rect 9419 14172 9483 14176
rect 9419 14116 9423 14172
rect 9423 14116 9479 14172
rect 9479 14116 9483 14172
rect 9419 14112 9483 14116
rect 9499 14172 9563 14176
rect 9499 14116 9503 14172
rect 9503 14116 9559 14172
rect 9559 14116 9563 14172
rect 9499 14112 9563 14116
rect 12318 14172 12382 14176
rect 12318 14116 12322 14172
rect 12322 14116 12378 14172
rect 12378 14116 12382 14172
rect 12318 14112 12382 14116
rect 12398 14172 12462 14176
rect 12398 14116 12402 14172
rect 12402 14116 12458 14172
rect 12458 14116 12462 14172
rect 12398 14112 12462 14116
rect 12478 14172 12542 14176
rect 12478 14116 12482 14172
rect 12482 14116 12538 14172
rect 12538 14116 12542 14172
rect 12478 14112 12542 14116
rect 12558 14172 12622 14176
rect 12558 14116 12562 14172
rect 12562 14116 12618 14172
rect 12618 14116 12622 14172
rect 12558 14112 12622 14116
rect 2481 13628 2545 13632
rect 2481 13572 2485 13628
rect 2485 13572 2541 13628
rect 2541 13572 2545 13628
rect 2481 13568 2545 13572
rect 2561 13628 2625 13632
rect 2561 13572 2565 13628
rect 2565 13572 2621 13628
rect 2621 13572 2625 13628
rect 2561 13568 2625 13572
rect 2641 13628 2705 13632
rect 2641 13572 2645 13628
rect 2645 13572 2701 13628
rect 2701 13572 2705 13628
rect 2641 13568 2705 13572
rect 2721 13628 2785 13632
rect 2721 13572 2725 13628
rect 2725 13572 2781 13628
rect 2781 13572 2785 13628
rect 2721 13568 2785 13572
rect 5540 13628 5604 13632
rect 5540 13572 5544 13628
rect 5544 13572 5600 13628
rect 5600 13572 5604 13628
rect 5540 13568 5604 13572
rect 5620 13628 5684 13632
rect 5620 13572 5624 13628
rect 5624 13572 5680 13628
rect 5680 13572 5684 13628
rect 5620 13568 5684 13572
rect 5700 13628 5764 13632
rect 5700 13572 5704 13628
rect 5704 13572 5760 13628
rect 5760 13572 5764 13628
rect 5700 13568 5764 13572
rect 5780 13628 5844 13632
rect 5780 13572 5784 13628
rect 5784 13572 5840 13628
rect 5840 13572 5844 13628
rect 5780 13568 5844 13572
rect 8599 13628 8663 13632
rect 8599 13572 8603 13628
rect 8603 13572 8659 13628
rect 8659 13572 8663 13628
rect 8599 13568 8663 13572
rect 8679 13628 8743 13632
rect 8679 13572 8683 13628
rect 8683 13572 8739 13628
rect 8739 13572 8743 13628
rect 8679 13568 8743 13572
rect 8759 13628 8823 13632
rect 8759 13572 8763 13628
rect 8763 13572 8819 13628
rect 8819 13572 8823 13628
rect 8759 13568 8823 13572
rect 8839 13628 8903 13632
rect 8839 13572 8843 13628
rect 8843 13572 8899 13628
rect 8899 13572 8903 13628
rect 8839 13568 8903 13572
rect 11658 13628 11722 13632
rect 11658 13572 11662 13628
rect 11662 13572 11718 13628
rect 11718 13572 11722 13628
rect 11658 13568 11722 13572
rect 11738 13628 11802 13632
rect 11738 13572 11742 13628
rect 11742 13572 11798 13628
rect 11798 13572 11802 13628
rect 11738 13568 11802 13572
rect 11818 13628 11882 13632
rect 11818 13572 11822 13628
rect 11822 13572 11878 13628
rect 11878 13572 11882 13628
rect 11818 13568 11882 13572
rect 11898 13628 11962 13632
rect 11898 13572 11902 13628
rect 11902 13572 11958 13628
rect 11958 13572 11962 13628
rect 11898 13568 11962 13572
rect 3141 13084 3205 13088
rect 3141 13028 3145 13084
rect 3145 13028 3201 13084
rect 3201 13028 3205 13084
rect 3141 13024 3205 13028
rect 3221 13084 3285 13088
rect 3221 13028 3225 13084
rect 3225 13028 3281 13084
rect 3281 13028 3285 13084
rect 3221 13024 3285 13028
rect 3301 13084 3365 13088
rect 3301 13028 3305 13084
rect 3305 13028 3361 13084
rect 3361 13028 3365 13084
rect 3301 13024 3365 13028
rect 3381 13084 3445 13088
rect 3381 13028 3385 13084
rect 3385 13028 3441 13084
rect 3441 13028 3445 13084
rect 3381 13024 3445 13028
rect 6200 13084 6264 13088
rect 6200 13028 6204 13084
rect 6204 13028 6260 13084
rect 6260 13028 6264 13084
rect 6200 13024 6264 13028
rect 6280 13084 6344 13088
rect 6280 13028 6284 13084
rect 6284 13028 6340 13084
rect 6340 13028 6344 13084
rect 6280 13024 6344 13028
rect 6360 13084 6424 13088
rect 6360 13028 6364 13084
rect 6364 13028 6420 13084
rect 6420 13028 6424 13084
rect 6360 13024 6424 13028
rect 6440 13084 6504 13088
rect 6440 13028 6444 13084
rect 6444 13028 6500 13084
rect 6500 13028 6504 13084
rect 6440 13024 6504 13028
rect 9259 13084 9323 13088
rect 9259 13028 9263 13084
rect 9263 13028 9319 13084
rect 9319 13028 9323 13084
rect 9259 13024 9323 13028
rect 9339 13084 9403 13088
rect 9339 13028 9343 13084
rect 9343 13028 9399 13084
rect 9399 13028 9403 13084
rect 9339 13024 9403 13028
rect 9419 13084 9483 13088
rect 9419 13028 9423 13084
rect 9423 13028 9479 13084
rect 9479 13028 9483 13084
rect 9419 13024 9483 13028
rect 9499 13084 9563 13088
rect 9499 13028 9503 13084
rect 9503 13028 9559 13084
rect 9559 13028 9563 13084
rect 9499 13024 9563 13028
rect 12318 13084 12382 13088
rect 12318 13028 12322 13084
rect 12322 13028 12378 13084
rect 12378 13028 12382 13084
rect 12318 13024 12382 13028
rect 12398 13084 12462 13088
rect 12398 13028 12402 13084
rect 12402 13028 12458 13084
rect 12458 13028 12462 13084
rect 12398 13024 12462 13028
rect 12478 13084 12542 13088
rect 12478 13028 12482 13084
rect 12482 13028 12538 13084
rect 12538 13028 12542 13084
rect 12478 13024 12542 13028
rect 12558 13084 12622 13088
rect 12558 13028 12562 13084
rect 12562 13028 12618 13084
rect 12618 13028 12622 13084
rect 12558 13024 12622 13028
rect 2481 12540 2545 12544
rect 2481 12484 2485 12540
rect 2485 12484 2541 12540
rect 2541 12484 2545 12540
rect 2481 12480 2545 12484
rect 2561 12540 2625 12544
rect 2561 12484 2565 12540
rect 2565 12484 2621 12540
rect 2621 12484 2625 12540
rect 2561 12480 2625 12484
rect 2641 12540 2705 12544
rect 2641 12484 2645 12540
rect 2645 12484 2701 12540
rect 2701 12484 2705 12540
rect 2641 12480 2705 12484
rect 2721 12540 2785 12544
rect 2721 12484 2725 12540
rect 2725 12484 2781 12540
rect 2781 12484 2785 12540
rect 2721 12480 2785 12484
rect 5540 12540 5604 12544
rect 5540 12484 5544 12540
rect 5544 12484 5600 12540
rect 5600 12484 5604 12540
rect 5540 12480 5604 12484
rect 5620 12540 5684 12544
rect 5620 12484 5624 12540
rect 5624 12484 5680 12540
rect 5680 12484 5684 12540
rect 5620 12480 5684 12484
rect 5700 12540 5764 12544
rect 5700 12484 5704 12540
rect 5704 12484 5760 12540
rect 5760 12484 5764 12540
rect 5700 12480 5764 12484
rect 5780 12540 5844 12544
rect 5780 12484 5784 12540
rect 5784 12484 5840 12540
rect 5840 12484 5844 12540
rect 5780 12480 5844 12484
rect 8599 12540 8663 12544
rect 8599 12484 8603 12540
rect 8603 12484 8659 12540
rect 8659 12484 8663 12540
rect 8599 12480 8663 12484
rect 8679 12540 8743 12544
rect 8679 12484 8683 12540
rect 8683 12484 8739 12540
rect 8739 12484 8743 12540
rect 8679 12480 8743 12484
rect 8759 12540 8823 12544
rect 8759 12484 8763 12540
rect 8763 12484 8819 12540
rect 8819 12484 8823 12540
rect 8759 12480 8823 12484
rect 8839 12540 8903 12544
rect 8839 12484 8843 12540
rect 8843 12484 8899 12540
rect 8899 12484 8903 12540
rect 8839 12480 8903 12484
rect 11658 12540 11722 12544
rect 11658 12484 11662 12540
rect 11662 12484 11718 12540
rect 11718 12484 11722 12540
rect 11658 12480 11722 12484
rect 11738 12540 11802 12544
rect 11738 12484 11742 12540
rect 11742 12484 11798 12540
rect 11798 12484 11802 12540
rect 11738 12480 11802 12484
rect 11818 12540 11882 12544
rect 11818 12484 11822 12540
rect 11822 12484 11878 12540
rect 11878 12484 11882 12540
rect 11818 12480 11882 12484
rect 11898 12540 11962 12544
rect 11898 12484 11902 12540
rect 11902 12484 11958 12540
rect 11958 12484 11962 12540
rect 11898 12480 11962 12484
rect 3141 11996 3205 12000
rect 3141 11940 3145 11996
rect 3145 11940 3201 11996
rect 3201 11940 3205 11996
rect 3141 11936 3205 11940
rect 3221 11996 3285 12000
rect 3221 11940 3225 11996
rect 3225 11940 3281 11996
rect 3281 11940 3285 11996
rect 3221 11936 3285 11940
rect 3301 11996 3365 12000
rect 3301 11940 3305 11996
rect 3305 11940 3361 11996
rect 3361 11940 3365 11996
rect 3301 11936 3365 11940
rect 3381 11996 3445 12000
rect 3381 11940 3385 11996
rect 3385 11940 3441 11996
rect 3441 11940 3445 11996
rect 3381 11936 3445 11940
rect 6200 11996 6264 12000
rect 6200 11940 6204 11996
rect 6204 11940 6260 11996
rect 6260 11940 6264 11996
rect 6200 11936 6264 11940
rect 6280 11996 6344 12000
rect 6280 11940 6284 11996
rect 6284 11940 6340 11996
rect 6340 11940 6344 11996
rect 6280 11936 6344 11940
rect 6360 11996 6424 12000
rect 6360 11940 6364 11996
rect 6364 11940 6420 11996
rect 6420 11940 6424 11996
rect 6360 11936 6424 11940
rect 6440 11996 6504 12000
rect 6440 11940 6444 11996
rect 6444 11940 6500 11996
rect 6500 11940 6504 11996
rect 6440 11936 6504 11940
rect 9259 11996 9323 12000
rect 9259 11940 9263 11996
rect 9263 11940 9319 11996
rect 9319 11940 9323 11996
rect 9259 11936 9323 11940
rect 9339 11996 9403 12000
rect 9339 11940 9343 11996
rect 9343 11940 9399 11996
rect 9399 11940 9403 11996
rect 9339 11936 9403 11940
rect 9419 11996 9483 12000
rect 9419 11940 9423 11996
rect 9423 11940 9479 11996
rect 9479 11940 9483 11996
rect 9419 11936 9483 11940
rect 9499 11996 9563 12000
rect 9499 11940 9503 11996
rect 9503 11940 9559 11996
rect 9559 11940 9563 11996
rect 9499 11936 9563 11940
rect 12318 11996 12382 12000
rect 12318 11940 12322 11996
rect 12322 11940 12378 11996
rect 12378 11940 12382 11996
rect 12318 11936 12382 11940
rect 12398 11996 12462 12000
rect 12398 11940 12402 11996
rect 12402 11940 12458 11996
rect 12458 11940 12462 11996
rect 12398 11936 12462 11940
rect 12478 11996 12542 12000
rect 12478 11940 12482 11996
rect 12482 11940 12538 11996
rect 12538 11940 12542 11996
rect 12478 11936 12542 11940
rect 12558 11996 12622 12000
rect 12558 11940 12562 11996
rect 12562 11940 12618 11996
rect 12618 11940 12622 11996
rect 12558 11936 12622 11940
rect 2481 11452 2545 11456
rect 2481 11396 2485 11452
rect 2485 11396 2541 11452
rect 2541 11396 2545 11452
rect 2481 11392 2545 11396
rect 2561 11452 2625 11456
rect 2561 11396 2565 11452
rect 2565 11396 2621 11452
rect 2621 11396 2625 11452
rect 2561 11392 2625 11396
rect 2641 11452 2705 11456
rect 2641 11396 2645 11452
rect 2645 11396 2701 11452
rect 2701 11396 2705 11452
rect 2641 11392 2705 11396
rect 2721 11452 2785 11456
rect 2721 11396 2725 11452
rect 2725 11396 2781 11452
rect 2781 11396 2785 11452
rect 2721 11392 2785 11396
rect 5540 11452 5604 11456
rect 5540 11396 5544 11452
rect 5544 11396 5600 11452
rect 5600 11396 5604 11452
rect 5540 11392 5604 11396
rect 5620 11452 5684 11456
rect 5620 11396 5624 11452
rect 5624 11396 5680 11452
rect 5680 11396 5684 11452
rect 5620 11392 5684 11396
rect 5700 11452 5764 11456
rect 5700 11396 5704 11452
rect 5704 11396 5760 11452
rect 5760 11396 5764 11452
rect 5700 11392 5764 11396
rect 5780 11452 5844 11456
rect 5780 11396 5784 11452
rect 5784 11396 5840 11452
rect 5840 11396 5844 11452
rect 5780 11392 5844 11396
rect 8599 11452 8663 11456
rect 8599 11396 8603 11452
rect 8603 11396 8659 11452
rect 8659 11396 8663 11452
rect 8599 11392 8663 11396
rect 8679 11452 8743 11456
rect 8679 11396 8683 11452
rect 8683 11396 8739 11452
rect 8739 11396 8743 11452
rect 8679 11392 8743 11396
rect 8759 11452 8823 11456
rect 8759 11396 8763 11452
rect 8763 11396 8819 11452
rect 8819 11396 8823 11452
rect 8759 11392 8823 11396
rect 8839 11452 8903 11456
rect 8839 11396 8843 11452
rect 8843 11396 8899 11452
rect 8899 11396 8903 11452
rect 8839 11392 8903 11396
rect 11658 11452 11722 11456
rect 11658 11396 11662 11452
rect 11662 11396 11718 11452
rect 11718 11396 11722 11452
rect 11658 11392 11722 11396
rect 11738 11452 11802 11456
rect 11738 11396 11742 11452
rect 11742 11396 11798 11452
rect 11798 11396 11802 11452
rect 11738 11392 11802 11396
rect 11818 11452 11882 11456
rect 11818 11396 11822 11452
rect 11822 11396 11878 11452
rect 11878 11396 11882 11452
rect 11818 11392 11882 11396
rect 11898 11452 11962 11456
rect 11898 11396 11902 11452
rect 11902 11396 11958 11452
rect 11958 11396 11962 11452
rect 11898 11392 11962 11396
rect 3141 10908 3205 10912
rect 3141 10852 3145 10908
rect 3145 10852 3201 10908
rect 3201 10852 3205 10908
rect 3141 10848 3205 10852
rect 3221 10908 3285 10912
rect 3221 10852 3225 10908
rect 3225 10852 3281 10908
rect 3281 10852 3285 10908
rect 3221 10848 3285 10852
rect 3301 10908 3365 10912
rect 3301 10852 3305 10908
rect 3305 10852 3361 10908
rect 3361 10852 3365 10908
rect 3301 10848 3365 10852
rect 3381 10908 3445 10912
rect 3381 10852 3385 10908
rect 3385 10852 3441 10908
rect 3441 10852 3445 10908
rect 3381 10848 3445 10852
rect 6200 10908 6264 10912
rect 6200 10852 6204 10908
rect 6204 10852 6260 10908
rect 6260 10852 6264 10908
rect 6200 10848 6264 10852
rect 6280 10908 6344 10912
rect 6280 10852 6284 10908
rect 6284 10852 6340 10908
rect 6340 10852 6344 10908
rect 6280 10848 6344 10852
rect 6360 10908 6424 10912
rect 6360 10852 6364 10908
rect 6364 10852 6420 10908
rect 6420 10852 6424 10908
rect 6360 10848 6424 10852
rect 6440 10908 6504 10912
rect 6440 10852 6444 10908
rect 6444 10852 6500 10908
rect 6500 10852 6504 10908
rect 6440 10848 6504 10852
rect 9259 10908 9323 10912
rect 9259 10852 9263 10908
rect 9263 10852 9319 10908
rect 9319 10852 9323 10908
rect 9259 10848 9323 10852
rect 9339 10908 9403 10912
rect 9339 10852 9343 10908
rect 9343 10852 9399 10908
rect 9399 10852 9403 10908
rect 9339 10848 9403 10852
rect 9419 10908 9483 10912
rect 9419 10852 9423 10908
rect 9423 10852 9479 10908
rect 9479 10852 9483 10908
rect 9419 10848 9483 10852
rect 9499 10908 9563 10912
rect 9499 10852 9503 10908
rect 9503 10852 9559 10908
rect 9559 10852 9563 10908
rect 9499 10848 9563 10852
rect 12318 10908 12382 10912
rect 12318 10852 12322 10908
rect 12322 10852 12378 10908
rect 12378 10852 12382 10908
rect 12318 10848 12382 10852
rect 12398 10908 12462 10912
rect 12398 10852 12402 10908
rect 12402 10852 12458 10908
rect 12458 10852 12462 10908
rect 12398 10848 12462 10852
rect 12478 10908 12542 10912
rect 12478 10852 12482 10908
rect 12482 10852 12538 10908
rect 12538 10852 12542 10908
rect 12478 10848 12542 10852
rect 12558 10908 12622 10912
rect 12558 10852 12562 10908
rect 12562 10852 12618 10908
rect 12618 10852 12622 10908
rect 12558 10848 12622 10852
rect 2481 10364 2545 10368
rect 2481 10308 2485 10364
rect 2485 10308 2541 10364
rect 2541 10308 2545 10364
rect 2481 10304 2545 10308
rect 2561 10364 2625 10368
rect 2561 10308 2565 10364
rect 2565 10308 2621 10364
rect 2621 10308 2625 10364
rect 2561 10304 2625 10308
rect 2641 10364 2705 10368
rect 2641 10308 2645 10364
rect 2645 10308 2701 10364
rect 2701 10308 2705 10364
rect 2641 10304 2705 10308
rect 2721 10364 2785 10368
rect 2721 10308 2725 10364
rect 2725 10308 2781 10364
rect 2781 10308 2785 10364
rect 2721 10304 2785 10308
rect 5540 10364 5604 10368
rect 5540 10308 5544 10364
rect 5544 10308 5600 10364
rect 5600 10308 5604 10364
rect 5540 10304 5604 10308
rect 5620 10364 5684 10368
rect 5620 10308 5624 10364
rect 5624 10308 5680 10364
rect 5680 10308 5684 10364
rect 5620 10304 5684 10308
rect 5700 10364 5764 10368
rect 5700 10308 5704 10364
rect 5704 10308 5760 10364
rect 5760 10308 5764 10364
rect 5700 10304 5764 10308
rect 5780 10364 5844 10368
rect 5780 10308 5784 10364
rect 5784 10308 5840 10364
rect 5840 10308 5844 10364
rect 5780 10304 5844 10308
rect 8599 10364 8663 10368
rect 8599 10308 8603 10364
rect 8603 10308 8659 10364
rect 8659 10308 8663 10364
rect 8599 10304 8663 10308
rect 8679 10364 8743 10368
rect 8679 10308 8683 10364
rect 8683 10308 8739 10364
rect 8739 10308 8743 10364
rect 8679 10304 8743 10308
rect 8759 10364 8823 10368
rect 8759 10308 8763 10364
rect 8763 10308 8819 10364
rect 8819 10308 8823 10364
rect 8759 10304 8823 10308
rect 8839 10364 8903 10368
rect 8839 10308 8843 10364
rect 8843 10308 8899 10364
rect 8899 10308 8903 10364
rect 8839 10304 8903 10308
rect 11658 10364 11722 10368
rect 11658 10308 11662 10364
rect 11662 10308 11718 10364
rect 11718 10308 11722 10364
rect 11658 10304 11722 10308
rect 11738 10364 11802 10368
rect 11738 10308 11742 10364
rect 11742 10308 11798 10364
rect 11798 10308 11802 10364
rect 11738 10304 11802 10308
rect 11818 10364 11882 10368
rect 11818 10308 11822 10364
rect 11822 10308 11878 10364
rect 11878 10308 11882 10364
rect 11818 10304 11882 10308
rect 11898 10364 11962 10368
rect 11898 10308 11902 10364
rect 11902 10308 11958 10364
rect 11958 10308 11962 10364
rect 11898 10304 11962 10308
rect 3141 9820 3205 9824
rect 3141 9764 3145 9820
rect 3145 9764 3201 9820
rect 3201 9764 3205 9820
rect 3141 9760 3205 9764
rect 3221 9820 3285 9824
rect 3221 9764 3225 9820
rect 3225 9764 3281 9820
rect 3281 9764 3285 9820
rect 3221 9760 3285 9764
rect 3301 9820 3365 9824
rect 3301 9764 3305 9820
rect 3305 9764 3361 9820
rect 3361 9764 3365 9820
rect 3301 9760 3365 9764
rect 3381 9820 3445 9824
rect 3381 9764 3385 9820
rect 3385 9764 3441 9820
rect 3441 9764 3445 9820
rect 3381 9760 3445 9764
rect 6200 9820 6264 9824
rect 6200 9764 6204 9820
rect 6204 9764 6260 9820
rect 6260 9764 6264 9820
rect 6200 9760 6264 9764
rect 6280 9820 6344 9824
rect 6280 9764 6284 9820
rect 6284 9764 6340 9820
rect 6340 9764 6344 9820
rect 6280 9760 6344 9764
rect 6360 9820 6424 9824
rect 6360 9764 6364 9820
rect 6364 9764 6420 9820
rect 6420 9764 6424 9820
rect 6360 9760 6424 9764
rect 6440 9820 6504 9824
rect 6440 9764 6444 9820
rect 6444 9764 6500 9820
rect 6500 9764 6504 9820
rect 6440 9760 6504 9764
rect 9259 9820 9323 9824
rect 9259 9764 9263 9820
rect 9263 9764 9319 9820
rect 9319 9764 9323 9820
rect 9259 9760 9323 9764
rect 9339 9820 9403 9824
rect 9339 9764 9343 9820
rect 9343 9764 9399 9820
rect 9399 9764 9403 9820
rect 9339 9760 9403 9764
rect 9419 9820 9483 9824
rect 9419 9764 9423 9820
rect 9423 9764 9479 9820
rect 9479 9764 9483 9820
rect 9419 9760 9483 9764
rect 9499 9820 9563 9824
rect 9499 9764 9503 9820
rect 9503 9764 9559 9820
rect 9559 9764 9563 9820
rect 9499 9760 9563 9764
rect 12318 9820 12382 9824
rect 12318 9764 12322 9820
rect 12322 9764 12378 9820
rect 12378 9764 12382 9820
rect 12318 9760 12382 9764
rect 12398 9820 12462 9824
rect 12398 9764 12402 9820
rect 12402 9764 12458 9820
rect 12458 9764 12462 9820
rect 12398 9760 12462 9764
rect 12478 9820 12542 9824
rect 12478 9764 12482 9820
rect 12482 9764 12538 9820
rect 12538 9764 12542 9820
rect 12478 9760 12542 9764
rect 12558 9820 12622 9824
rect 12558 9764 12562 9820
rect 12562 9764 12618 9820
rect 12618 9764 12622 9820
rect 12558 9760 12622 9764
rect 2481 9276 2545 9280
rect 2481 9220 2485 9276
rect 2485 9220 2541 9276
rect 2541 9220 2545 9276
rect 2481 9216 2545 9220
rect 2561 9276 2625 9280
rect 2561 9220 2565 9276
rect 2565 9220 2621 9276
rect 2621 9220 2625 9276
rect 2561 9216 2625 9220
rect 2641 9276 2705 9280
rect 2641 9220 2645 9276
rect 2645 9220 2701 9276
rect 2701 9220 2705 9276
rect 2641 9216 2705 9220
rect 2721 9276 2785 9280
rect 2721 9220 2725 9276
rect 2725 9220 2781 9276
rect 2781 9220 2785 9276
rect 2721 9216 2785 9220
rect 5540 9276 5604 9280
rect 5540 9220 5544 9276
rect 5544 9220 5600 9276
rect 5600 9220 5604 9276
rect 5540 9216 5604 9220
rect 5620 9276 5684 9280
rect 5620 9220 5624 9276
rect 5624 9220 5680 9276
rect 5680 9220 5684 9276
rect 5620 9216 5684 9220
rect 5700 9276 5764 9280
rect 5700 9220 5704 9276
rect 5704 9220 5760 9276
rect 5760 9220 5764 9276
rect 5700 9216 5764 9220
rect 5780 9276 5844 9280
rect 5780 9220 5784 9276
rect 5784 9220 5840 9276
rect 5840 9220 5844 9276
rect 5780 9216 5844 9220
rect 8599 9276 8663 9280
rect 8599 9220 8603 9276
rect 8603 9220 8659 9276
rect 8659 9220 8663 9276
rect 8599 9216 8663 9220
rect 8679 9276 8743 9280
rect 8679 9220 8683 9276
rect 8683 9220 8739 9276
rect 8739 9220 8743 9276
rect 8679 9216 8743 9220
rect 8759 9276 8823 9280
rect 8759 9220 8763 9276
rect 8763 9220 8819 9276
rect 8819 9220 8823 9276
rect 8759 9216 8823 9220
rect 8839 9276 8903 9280
rect 8839 9220 8843 9276
rect 8843 9220 8899 9276
rect 8899 9220 8903 9276
rect 8839 9216 8903 9220
rect 11658 9276 11722 9280
rect 11658 9220 11662 9276
rect 11662 9220 11718 9276
rect 11718 9220 11722 9276
rect 11658 9216 11722 9220
rect 11738 9276 11802 9280
rect 11738 9220 11742 9276
rect 11742 9220 11798 9276
rect 11798 9220 11802 9276
rect 11738 9216 11802 9220
rect 11818 9276 11882 9280
rect 11818 9220 11822 9276
rect 11822 9220 11878 9276
rect 11878 9220 11882 9276
rect 11818 9216 11882 9220
rect 11898 9276 11962 9280
rect 11898 9220 11902 9276
rect 11902 9220 11958 9276
rect 11958 9220 11962 9276
rect 11898 9216 11962 9220
rect 3141 8732 3205 8736
rect 3141 8676 3145 8732
rect 3145 8676 3201 8732
rect 3201 8676 3205 8732
rect 3141 8672 3205 8676
rect 3221 8732 3285 8736
rect 3221 8676 3225 8732
rect 3225 8676 3281 8732
rect 3281 8676 3285 8732
rect 3221 8672 3285 8676
rect 3301 8732 3365 8736
rect 3301 8676 3305 8732
rect 3305 8676 3361 8732
rect 3361 8676 3365 8732
rect 3301 8672 3365 8676
rect 3381 8732 3445 8736
rect 3381 8676 3385 8732
rect 3385 8676 3441 8732
rect 3441 8676 3445 8732
rect 3381 8672 3445 8676
rect 6200 8732 6264 8736
rect 6200 8676 6204 8732
rect 6204 8676 6260 8732
rect 6260 8676 6264 8732
rect 6200 8672 6264 8676
rect 6280 8732 6344 8736
rect 6280 8676 6284 8732
rect 6284 8676 6340 8732
rect 6340 8676 6344 8732
rect 6280 8672 6344 8676
rect 6360 8732 6424 8736
rect 6360 8676 6364 8732
rect 6364 8676 6420 8732
rect 6420 8676 6424 8732
rect 6360 8672 6424 8676
rect 6440 8732 6504 8736
rect 6440 8676 6444 8732
rect 6444 8676 6500 8732
rect 6500 8676 6504 8732
rect 6440 8672 6504 8676
rect 9259 8732 9323 8736
rect 9259 8676 9263 8732
rect 9263 8676 9319 8732
rect 9319 8676 9323 8732
rect 9259 8672 9323 8676
rect 9339 8732 9403 8736
rect 9339 8676 9343 8732
rect 9343 8676 9399 8732
rect 9399 8676 9403 8732
rect 9339 8672 9403 8676
rect 9419 8732 9483 8736
rect 9419 8676 9423 8732
rect 9423 8676 9479 8732
rect 9479 8676 9483 8732
rect 9419 8672 9483 8676
rect 9499 8732 9563 8736
rect 9499 8676 9503 8732
rect 9503 8676 9559 8732
rect 9559 8676 9563 8732
rect 9499 8672 9563 8676
rect 12318 8732 12382 8736
rect 12318 8676 12322 8732
rect 12322 8676 12378 8732
rect 12378 8676 12382 8732
rect 12318 8672 12382 8676
rect 12398 8732 12462 8736
rect 12398 8676 12402 8732
rect 12402 8676 12458 8732
rect 12458 8676 12462 8732
rect 12398 8672 12462 8676
rect 12478 8732 12542 8736
rect 12478 8676 12482 8732
rect 12482 8676 12538 8732
rect 12538 8676 12542 8732
rect 12478 8672 12542 8676
rect 12558 8732 12622 8736
rect 12558 8676 12562 8732
rect 12562 8676 12618 8732
rect 12618 8676 12622 8732
rect 12558 8672 12622 8676
rect 2481 8188 2545 8192
rect 2481 8132 2485 8188
rect 2485 8132 2541 8188
rect 2541 8132 2545 8188
rect 2481 8128 2545 8132
rect 2561 8188 2625 8192
rect 2561 8132 2565 8188
rect 2565 8132 2621 8188
rect 2621 8132 2625 8188
rect 2561 8128 2625 8132
rect 2641 8188 2705 8192
rect 2641 8132 2645 8188
rect 2645 8132 2701 8188
rect 2701 8132 2705 8188
rect 2641 8128 2705 8132
rect 2721 8188 2785 8192
rect 2721 8132 2725 8188
rect 2725 8132 2781 8188
rect 2781 8132 2785 8188
rect 2721 8128 2785 8132
rect 5540 8188 5604 8192
rect 5540 8132 5544 8188
rect 5544 8132 5600 8188
rect 5600 8132 5604 8188
rect 5540 8128 5604 8132
rect 5620 8188 5684 8192
rect 5620 8132 5624 8188
rect 5624 8132 5680 8188
rect 5680 8132 5684 8188
rect 5620 8128 5684 8132
rect 5700 8188 5764 8192
rect 5700 8132 5704 8188
rect 5704 8132 5760 8188
rect 5760 8132 5764 8188
rect 5700 8128 5764 8132
rect 5780 8188 5844 8192
rect 5780 8132 5784 8188
rect 5784 8132 5840 8188
rect 5840 8132 5844 8188
rect 5780 8128 5844 8132
rect 8599 8188 8663 8192
rect 8599 8132 8603 8188
rect 8603 8132 8659 8188
rect 8659 8132 8663 8188
rect 8599 8128 8663 8132
rect 8679 8188 8743 8192
rect 8679 8132 8683 8188
rect 8683 8132 8739 8188
rect 8739 8132 8743 8188
rect 8679 8128 8743 8132
rect 8759 8188 8823 8192
rect 8759 8132 8763 8188
rect 8763 8132 8819 8188
rect 8819 8132 8823 8188
rect 8759 8128 8823 8132
rect 8839 8188 8903 8192
rect 8839 8132 8843 8188
rect 8843 8132 8899 8188
rect 8899 8132 8903 8188
rect 8839 8128 8903 8132
rect 11658 8188 11722 8192
rect 11658 8132 11662 8188
rect 11662 8132 11718 8188
rect 11718 8132 11722 8188
rect 11658 8128 11722 8132
rect 11738 8188 11802 8192
rect 11738 8132 11742 8188
rect 11742 8132 11798 8188
rect 11798 8132 11802 8188
rect 11738 8128 11802 8132
rect 11818 8188 11882 8192
rect 11818 8132 11822 8188
rect 11822 8132 11878 8188
rect 11878 8132 11882 8188
rect 11818 8128 11882 8132
rect 11898 8188 11962 8192
rect 11898 8132 11902 8188
rect 11902 8132 11958 8188
rect 11958 8132 11962 8188
rect 11898 8128 11962 8132
rect 3141 7644 3205 7648
rect 3141 7588 3145 7644
rect 3145 7588 3201 7644
rect 3201 7588 3205 7644
rect 3141 7584 3205 7588
rect 3221 7644 3285 7648
rect 3221 7588 3225 7644
rect 3225 7588 3281 7644
rect 3281 7588 3285 7644
rect 3221 7584 3285 7588
rect 3301 7644 3365 7648
rect 3301 7588 3305 7644
rect 3305 7588 3361 7644
rect 3361 7588 3365 7644
rect 3301 7584 3365 7588
rect 3381 7644 3445 7648
rect 3381 7588 3385 7644
rect 3385 7588 3441 7644
rect 3441 7588 3445 7644
rect 3381 7584 3445 7588
rect 6200 7644 6264 7648
rect 6200 7588 6204 7644
rect 6204 7588 6260 7644
rect 6260 7588 6264 7644
rect 6200 7584 6264 7588
rect 6280 7644 6344 7648
rect 6280 7588 6284 7644
rect 6284 7588 6340 7644
rect 6340 7588 6344 7644
rect 6280 7584 6344 7588
rect 6360 7644 6424 7648
rect 6360 7588 6364 7644
rect 6364 7588 6420 7644
rect 6420 7588 6424 7644
rect 6360 7584 6424 7588
rect 6440 7644 6504 7648
rect 6440 7588 6444 7644
rect 6444 7588 6500 7644
rect 6500 7588 6504 7644
rect 6440 7584 6504 7588
rect 9259 7644 9323 7648
rect 9259 7588 9263 7644
rect 9263 7588 9319 7644
rect 9319 7588 9323 7644
rect 9259 7584 9323 7588
rect 9339 7644 9403 7648
rect 9339 7588 9343 7644
rect 9343 7588 9399 7644
rect 9399 7588 9403 7644
rect 9339 7584 9403 7588
rect 9419 7644 9483 7648
rect 9419 7588 9423 7644
rect 9423 7588 9479 7644
rect 9479 7588 9483 7644
rect 9419 7584 9483 7588
rect 9499 7644 9563 7648
rect 9499 7588 9503 7644
rect 9503 7588 9559 7644
rect 9559 7588 9563 7644
rect 9499 7584 9563 7588
rect 12318 7644 12382 7648
rect 12318 7588 12322 7644
rect 12322 7588 12378 7644
rect 12378 7588 12382 7644
rect 12318 7584 12382 7588
rect 12398 7644 12462 7648
rect 12398 7588 12402 7644
rect 12402 7588 12458 7644
rect 12458 7588 12462 7644
rect 12398 7584 12462 7588
rect 12478 7644 12542 7648
rect 12478 7588 12482 7644
rect 12482 7588 12538 7644
rect 12538 7588 12542 7644
rect 12478 7584 12542 7588
rect 12558 7644 12622 7648
rect 12558 7588 12562 7644
rect 12562 7588 12618 7644
rect 12618 7588 12622 7644
rect 12558 7584 12622 7588
rect 2481 7100 2545 7104
rect 2481 7044 2485 7100
rect 2485 7044 2541 7100
rect 2541 7044 2545 7100
rect 2481 7040 2545 7044
rect 2561 7100 2625 7104
rect 2561 7044 2565 7100
rect 2565 7044 2621 7100
rect 2621 7044 2625 7100
rect 2561 7040 2625 7044
rect 2641 7100 2705 7104
rect 2641 7044 2645 7100
rect 2645 7044 2701 7100
rect 2701 7044 2705 7100
rect 2641 7040 2705 7044
rect 2721 7100 2785 7104
rect 2721 7044 2725 7100
rect 2725 7044 2781 7100
rect 2781 7044 2785 7100
rect 2721 7040 2785 7044
rect 5540 7100 5604 7104
rect 5540 7044 5544 7100
rect 5544 7044 5600 7100
rect 5600 7044 5604 7100
rect 5540 7040 5604 7044
rect 5620 7100 5684 7104
rect 5620 7044 5624 7100
rect 5624 7044 5680 7100
rect 5680 7044 5684 7100
rect 5620 7040 5684 7044
rect 5700 7100 5764 7104
rect 5700 7044 5704 7100
rect 5704 7044 5760 7100
rect 5760 7044 5764 7100
rect 5700 7040 5764 7044
rect 5780 7100 5844 7104
rect 5780 7044 5784 7100
rect 5784 7044 5840 7100
rect 5840 7044 5844 7100
rect 5780 7040 5844 7044
rect 8599 7100 8663 7104
rect 8599 7044 8603 7100
rect 8603 7044 8659 7100
rect 8659 7044 8663 7100
rect 8599 7040 8663 7044
rect 8679 7100 8743 7104
rect 8679 7044 8683 7100
rect 8683 7044 8739 7100
rect 8739 7044 8743 7100
rect 8679 7040 8743 7044
rect 8759 7100 8823 7104
rect 8759 7044 8763 7100
rect 8763 7044 8819 7100
rect 8819 7044 8823 7100
rect 8759 7040 8823 7044
rect 8839 7100 8903 7104
rect 8839 7044 8843 7100
rect 8843 7044 8899 7100
rect 8899 7044 8903 7100
rect 8839 7040 8903 7044
rect 11658 7100 11722 7104
rect 11658 7044 11662 7100
rect 11662 7044 11718 7100
rect 11718 7044 11722 7100
rect 11658 7040 11722 7044
rect 11738 7100 11802 7104
rect 11738 7044 11742 7100
rect 11742 7044 11798 7100
rect 11798 7044 11802 7100
rect 11738 7040 11802 7044
rect 11818 7100 11882 7104
rect 11818 7044 11822 7100
rect 11822 7044 11878 7100
rect 11878 7044 11882 7100
rect 11818 7040 11882 7044
rect 11898 7100 11962 7104
rect 11898 7044 11902 7100
rect 11902 7044 11958 7100
rect 11958 7044 11962 7100
rect 11898 7040 11962 7044
rect 3141 6556 3205 6560
rect 3141 6500 3145 6556
rect 3145 6500 3201 6556
rect 3201 6500 3205 6556
rect 3141 6496 3205 6500
rect 3221 6556 3285 6560
rect 3221 6500 3225 6556
rect 3225 6500 3281 6556
rect 3281 6500 3285 6556
rect 3221 6496 3285 6500
rect 3301 6556 3365 6560
rect 3301 6500 3305 6556
rect 3305 6500 3361 6556
rect 3361 6500 3365 6556
rect 3301 6496 3365 6500
rect 3381 6556 3445 6560
rect 3381 6500 3385 6556
rect 3385 6500 3441 6556
rect 3441 6500 3445 6556
rect 3381 6496 3445 6500
rect 6200 6556 6264 6560
rect 6200 6500 6204 6556
rect 6204 6500 6260 6556
rect 6260 6500 6264 6556
rect 6200 6496 6264 6500
rect 6280 6556 6344 6560
rect 6280 6500 6284 6556
rect 6284 6500 6340 6556
rect 6340 6500 6344 6556
rect 6280 6496 6344 6500
rect 6360 6556 6424 6560
rect 6360 6500 6364 6556
rect 6364 6500 6420 6556
rect 6420 6500 6424 6556
rect 6360 6496 6424 6500
rect 6440 6556 6504 6560
rect 6440 6500 6444 6556
rect 6444 6500 6500 6556
rect 6500 6500 6504 6556
rect 6440 6496 6504 6500
rect 9259 6556 9323 6560
rect 9259 6500 9263 6556
rect 9263 6500 9319 6556
rect 9319 6500 9323 6556
rect 9259 6496 9323 6500
rect 9339 6556 9403 6560
rect 9339 6500 9343 6556
rect 9343 6500 9399 6556
rect 9399 6500 9403 6556
rect 9339 6496 9403 6500
rect 9419 6556 9483 6560
rect 9419 6500 9423 6556
rect 9423 6500 9479 6556
rect 9479 6500 9483 6556
rect 9419 6496 9483 6500
rect 9499 6556 9563 6560
rect 9499 6500 9503 6556
rect 9503 6500 9559 6556
rect 9559 6500 9563 6556
rect 9499 6496 9563 6500
rect 12318 6556 12382 6560
rect 12318 6500 12322 6556
rect 12322 6500 12378 6556
rect 12378 6500 12382 6556
rect 12318 6496 12382 6500
rect 12398 6556 12462 6560
rect 12398 6500 12402 6556
rect 12402 6500 12458 6556
rect 12458 6500 12462 6556
rect 12398 6496 12462 6500
rect 12478 6556 12542 6560
rect 12478 6500 12482 6556
rect 12482 6500 12538 6556
rect 12538 6500 12542 6556
rect 12478 6496 12542 6500
rect 12558 6556 12622 6560
rect 12558 6500 12562 6556
rect 12562 6500 12618 6556
rect 12618 6500 12622 6556
rect 12558 6496 12622 6500
rect 2481 6012 2545 6016
rect 2481 5956 2485 6012
rect 2485 5956 2541 6012
rect 2541 5956 2545 6012
rect 2481 5952 2545 5956
rect 2561 6012 2625 6016
rect 2561 5956 2565 6012
rect 2565 5956 2621 6012
rect 2621 5956 2625 6012
rect 2561 5952 2625 5956
rect 2641 6012 2705 6016
rect 2641 5956 2645 6012
rect 2645 5956 2701 6012
rect 2701 5956 2705 6012
rect 2641 5952 2705 5956
rect 2721 6012 2785 6016
rect 2721 5956 2725 6012
rect 2725 5956 2781 6012
rect 2781 5956 2785 6012
rect 2721 5952 2785 5956
rect 5540 6012 5604 6016
rect 5540 5956 5544 6012
rect 5544 5956 5600 6012
rect 5600 5956 5604 6012
rect 5540 5952 5604 5956
rect 5620 6012 5684 6016
rect 5620 5956 5624 6012
rect 5624 5956 5680 6012
rect 5680 5956 5684 6012
rect 5620 5952 5684 5956
rect 5700 6012 5764 6016
rect 5700 5956 5704 6012
rect 5704 5956 5760 6012
rect 5760 5956 5764 6012
rect 5700 5952 5764 5956
rect 5780 6012 5844 6016
rect 5780 5956 5784 6012
rect 5784 5956 5840 6012
rect 5840 5956 5844 6012
rect 5780 5952 5844 5956
rect 8599 6012 8663 6016
rect 8599 5956 8603 6012
rect 8603 5956 8659 6012
rect 8659 5956 8663 6012
rect 8599 5952 8663 5956
rect 8679 6012 8743 6016
rect 8679 5956 8683 6012
rect 8683 5956 8739 6012
rect 8739 5956 8743 6012
rect 8679 5952 8743 5956
rect 8759 6012 8823 6016
rect 8759 5956 8763 6012
rect 8763 5956 8819 6012
rect 8819 5956 8823 6012
rect 8759 5952 8823 5956
rect 8839 6012 8903 6016
rect 8839 5956 8843 6012
rect 8843 5956 8899 6012
rect 8899 5956 8903 6012
rect 8839 5952 8903 5956
rect 11658 6012 11722 6016
rect 11658 5956 11662 6012
rect 11662 5956 11718 6012
rect 11718 5956 11722 6012
rect 11658 5952 11722 5956
rect 11738 6012 11802 6016
rect 11738 5956 11742 6012
rect 11742 5956 11798 6012
rect 11798 5956 11802 6012
rect 11738 5952 11802 5956
rect 11818 6012 11882 6016
rect 11818 5956 11822 6012
rect 11822 5956 11878 6012
rect 11878 5956 11882 6012
rect 11818 5952 11882 5956
rect 11898 6012 11962 6016
rect 11898 5956 11902 6012
rect 11902 5956 11958 6012
rect 11958 5956 11962 6012
rect 11898 5952 11962 5956
rect 3141 5468 3205 5472
rect 3141 5412 3145 5468
rect 3145 5412 3201 5468
rect 3201 5412 3205 5468
rect 3141 5408 3205 5412
rect 3221 5468 3285 5472
rect 3221 5412 3225 5468
rect 3225 5412 3281 5468
rect 3281 5412 3285 5468
rect 3221 5408 3285 5412
rect 3301 5468 3365 5472
rect 3301 5412 3305 5468
rect 3305 5412 3361 5468
rect 3361 5412 3365 5468
rect 3301 5408 3365 5412
rect 3381 5468 3445 5472
rect 3381 5412 3385 5468
rect 3385 5412 3441 5468
rect 3441 5412 3445 5468
rect 3381 5408 3445 5412
rect 6200 5468 6264 5472
rect 6200 5412 6204 5468
rect 6204 5412 6260 5468
rect 6260 5412 6264 5468
rect 6200 5408 6264 5412
rect 6280 5468 6344 5472
rect 6280 5412 6284 5468
rect 6284 5412 6340 5468
rect 6340 5412 6344 5468
rect 6280 5408 6344 5412
rect 6360 5468 6424 5472
rect 6360 5412 6364 5468
rect 6364 5412 6420 5468
rect 6420 5412 6424 5468
rect 6360 5408 6424 5412
rect 6440 5468 6504 5472
rect 6440 5412 6444 5468
rect 6444 5412 6500 5468
rect 6500 5412 6504 5468
rect 6440 5408 6504 5412
rect 9259 5468 9323 5472
rect 9259 5412 9263 5468
rect 9263 5412 9319 5468
rect 9319 5412 9323 5468
rect 9259 5408 9323 5412
rect 9339 5468 9403 5472
rect 9339 5412 9343 5468
rect 9343 5412 9399 5468
rect 9399 5412 9403 5468
rect 9339 5408 9403 5412
rect 9419 5468 9483 5472
rect 9419 5412 9423 5468
rect 9423 5412 9479 5468
rect 9479 5412 9483 5468
rect 9419 5408 9483 5412
rect 9499 5468 9563 5472
rect 9499 5412 9503 5468
rect 9503 5412 9559 5468
rect 9559 5412 9563 5468
rect 9499 5408 9563 5412
rect 12318 5468 12382 5472
rect 12318 5412 12322 5468
rect 12322 5412 12378 5468
rect 12378 5412 12382 5468
rect 12318 5408 12382 5412
rect 12398 5468 12462 5472
rect 12398 5412 12402 5468
rect 12402 5412 12458 5468
rect 12458 5412 12462 5468
rect 12398 5408 12462 5412
rect 12478 5468 12542 5472
rect 12478 5412 12482 5468
rect 12482 5412 12538 5468
rect 12538 5412 12542 5468
rect 12478 5408 12542 5412
rect 12558 5468 12622 5472
rect 12558 5412 12562 5468
rect 12562 5412 12618 5468
rect 12618 5412 12622 5468
rect 12558 5408 12622 5412
rect 2481 4924 2545 4928
rect 2481 4868 2485 4924
rect 2485 4868 2541 4924
rect 2541 4868 2545 4924
rect 2481 4864 2545 4868
rect 2561 4924 2625 4928
rect 2561 4868 2565 4924
rect 2565 4868 2621 4924
rect 2621 4868 2625 4924
rect 2561 4864 2625 4868
rect 2641 4924 2705 4928
rect 2641 4868 2645 4924
rect 2645 4868 2701 4924
rect 2701 4868 2705 4924
rect 2641 4864 2705 4868
rect 2721 4924 2785 4928
rect 2721 4868 2725 4924
rect 2725 4868 2781 4924
rect 2781 4868 2785 4924
rect 2721 4864 2785 4868
rect 5540 4924 5604 4928
rect 5540 4868 5544 4924
rect 5544 4868 5600 4924
rect 5600 4868 5604 4924
rect 5540 4864 5604 4868
rect 5620 4924 5684 4928
rect 5620 4868 5624 4924
rect 5624 4868 5680 4924
rect 5680 4868 5684 4924
rect 5620 4864 5684 4868
rect 5700 4924 5764 4928
rect 5700 4868 5704 4924
rect 5704 4868 5760 4924
rect 5760 4868 5764 4924
rect 5700 4864 5764 4868
rect 5780 4924 5844 4928
rect 5780 4868 5784 4924
rect 5784 4868 5840 4924
rect 5840 4868 5844 4924
rect 5780 4864 5844 4868
rect 8599 4924 8663 4928
rect 8599 4868 8603 4924
rect 8603 4868 8659 4924
rect 8659 4868 8663 4924
rect 8599 4864 8663 4868
rect 8679 4924 8743 4928
rect 8679 4868 8683 4924
rect 8683 4868 8739 4924
rect 8739 4868 8743 4924
rect 8679 4864 8743 4868
rect 8759 4924 8823 4928
rect 8759 4868 8763 4924
rect 8763 4868 8819 4924
rect 8819 4868 8823 4924
rect 8759 4864 8823 4868
rect 8839 4924 8903 4928
rect 8839 4868 8843 4924
rect 8843 4868 8899 4924
rect 8899 4868 8903 4924
rect 8839 4864 8903 4868
rect 11658 4924 11722 4928
rect 11658 4868 11662 4924
rect 11662 4868 11718 4924
rect 11718 4868 11722 4924
rect 11658 4864 11722 4868
rect 11738 4924 11802 4928
rect 11738 4868 11742 4924
rect 11742 4868 11798 4924
rect 11798 4868 11802 4924
rect 11738 4864 11802 4868
rect 11818 4924 11882 4928
rect 11818 4868 11822 4924
rect 11822 4868 11878 4924
rect 11878 4868 11882 4924
rect 11818 4864 11882 4868
rect 11898 4924 11962 4928
rect 11898 4868 11902 4924
rect 11902 4868 11958 4924
rect 11958 4868 11962 4924
rect 11898 4864 11962 4868
rect 3141 4380 3205 4384
rect 3141 4324 3145 4380
rect 3145 4324 3201 4380
rect 3201 4324 3205 4380
rect 3141 4320 3205 4324
rect 3221 4380 3285 4384
rect 3221 4324 3225 4380
rect 3225 4324 3281 4380
rect 3281 4324 3285 4380
rect 3221 4320 3285 4324
rect 3301 4380 3365 4384
rect 3301 4324 3305 4380
rect 3305 4324 3361 4380
rect 3361 4324 3365 4380
rect 3301 4320 3365 4324
rect 3381 4380 3445 4384
rect 3381 4324 3385 4380
rect 3385 4324 3441 4380
rect 3441 4324 3445 4380
rect 3381 4320 3445 4324
rect 6200 4380 6264 4384
rect 6200 4324 6204 4380
rect 6204 4324 6260 4380
rect 6260 4324 6264 4380
rect 6200 4320 6264 4324
rect 6280 4380 6344 4384
rect 6280 4324 6284 4380
rect 6284 4324 6340 4380
rect 6340 4324 6344 4380
rect 6280 4320 6344 4324
rect 6360 4380 6424 4384
rect 6360 4324 6364 4380
rect 6364 4324 6420 4380
rect 6420 4324 6424 4380
rect 6360 4320 6424 4324
rect 6440 4380 6504 4384
rect 6440 4324 6444 4380
rect 6444 4324 6500 4380
rect 6500 4324 6504 4380
rect 6440 4320 6504 4324
rect 9259 4380 9323 4384
rect 9259 4324 9263 4380
rect 9263 4324 9319 4380
rect 9319 4324 9323 4380
rect 9259 4320 9323 4324
rect 9339 4380 9403 4384
rect 9339 4324 9343 4380
rect 9343 4324 9399 4380
rect 9399 4324 9403 4380
rect 9339 4320 9403 4324
rect 9419 4380 9483 4384
rect 9419 4324 9423 4380
rect 9423 4324 9479 4380
rect 9479 4324 9483 4380
rect 9419 4320 9483 4324
rect 9499 4380 9563 4384
rect 9499 4324 9503 4380
rect 9503 4324 9559 4380
rect 9559 4324 9563 4380
rect 9499 4320 9563 4324
rect 12318 4380 12382 4384
rect 12318 4324 12322 4380
rect 12322 4324 12378 4380
rect 12378 4324 12382 4380
rect 12318 4320 12382 4324
rect 12398 4380 12462 4384
rect 12398 4324 12402 4380
rect 12402 4324 12458 4380
rect 12458 4324 12462 4380
rect 12398 4320 12462 4324
rect 12478 4380 12542 4384
rect 12478 4324 12482 4380
rect 12482 4324 12538 4380
rect 12538 4324 12542 4380
rect 12478 4320 12542 4324
rect 12558 4380 12622 4384
rect 12558 4324 12562 4380
rect 12562 4324 12618 4380
rect 12618 4324 12622 4380
rect 12558 4320 12622 4324
rect 2481 3836 2545 3840
rect 2481 3780 2485 3836
rect 2485 3780 2541 3836
rect 2541 3780 2545 3836
rect 2481 3776 2545 3780
rect 2561 3836 2625 3840
rect 2561 3780 2565 3836
rect 2565 3780 2621 3836
rect 2621 3780 2625 3836
rect 2561 3776 2625 3780
rect 2641 3836 2705 3840
rect 2641 3780 2645 3836
rect 2645 3780 2701 3836
rect 2701 3780 2705 3836
rect 2641 3776 2705 3780
rect 2721 3836 2785 3840
rect 2721 3780 2725 3836
rect 2725 3780 2781 3836
rect 2781 3780 2785 3836
rect 2721 3776 2785 3780
rect 5540 3836 5604 3840
rect 5540 3780 5544 3836
rect 5544 3780 5600 3836
rect 5600 3780 5604 3836
rect 5540 3776 5604 3780
rect 5620 3836 5684 3840
rect 5620 3780 5624 3836
rect 5624 3780 5680 3836
rect 5680 3780 5684 3836
rect 5620 3776 5684 3780
rect 5700 3836 5764 3840
rect 5700 3780 5704 3836
rect 5704 3780 5760 3836
rect 5760 3780 5764 3836
rect 5700 3776 5764 3780
rect 5780 3836 5844 3840
rect 5780 3780 5784 3836
rect 5784 3780 5840 3836
rect 5840 3780 5844 3836
rect 5780 3776 5844 3780
rect 8599 3836 8663 3840
rect 8599 3780 8603 3836
rect 8603 3780 8659 3836
rect 8659 3780 8663 3836
rect 8599 3776 8663 3780
rect 8679 3836 8743 3840
rect 8679 3780 8683 3836
rect 8683 3780 8739 3836
rect 8739 3780 8743 3836
rect 8679 3776 8743 3780
rect 8759 3836 8823 3840
rect 8759 3780 8763 3836
rect 8763 3780 8819 3836
rect 8819 3780 8823 3836
rect 8759 3776 8823 3780
rect 8839 3836 8903 3840
rect 8839 3780 8843 3836
rect 8843 3780 8899 3836
rect 8899 3780 8903 3836
rect 8839 3776 8903 3780
rect 11658 3836 11722 3840
rect 11658 3780 11662 3836
rect 11662 3780 11718 3836
rect 11718 3780 11722 3836
rect 11658 3776 11722 3780
rect 11738 3836 11802 3840
rect 11738 3780 11742 3836
rect 11742 3780 11798 3836
rect 11798 3780 11802 3836
rect 11738 3776 11802 3780
rect 11818 3836 11882 3840
rect 11818 3780 11822 3836
rect 11822 3780 11878 3836
rect 11878 3780 11882 3836
rect 11818 3776 11882 3780
rect 11898 3836 11962 3840
rect 11898 3780 11902 3836
rect 11902 3780 11958 3836
rect 11958 3780 11962 3836
rect 11898 3776 11962 3780
rect 3141 3292 3205 3296
rect 3141 3236 3145 3292
rect 3145 3236 3201 3292
rect 3201 3236 3205 3292
rect 3141 3232 3205 3236
rect 3221 3292 3285 3296
rect 3221 3236 3225 3292
rect 3225 3236 3281 3292
rect 3281 3236 3285 3292
rect 3221 3232 3285 3236
rect 3301 3292 3365 3296
rect 3301 3236 3305 3292
rect 3305 3236 3361 3292
rect 3361 3236 3365 3292
rect 3301 3232 3365 3236
rect 3381 3292 3445 3296
rect 3381 3236 3385 3292
rect 3385 3236 3441 3292
rect 3441 3236 3445 3292
rect 3381 3232 3445 3236
rect 6200 3292 6264 3296
rect 6200 3236 6204 3292
rect 6204 3236 6260 3292
rect 6260 3236 6264 3292
rect 6200 3232 6264 3236
rect 6280 3292 6344 3296
rect 6280 3236 6284 3292
rect 6284 3236 6340 3292
rect 6340 3236 6344 3292
rect 6280 3232 6344 3236
rect 6360 3292 6424 3296
rect 6360 3236 6364 3292
rect 6364 3236 6420 3292
rect 6420 3236 6424 3292
rect 6360 3232 6424 3236
rect 6440 3292 6504 3296
rect 6440 3236 6444 3292
rect 6444 3236 6500 3292
rect 6500 3236 6504 3292
rect 6440 3232 6504 3236
rect 9259 3292 9323 3296
rect 9259 3236 9263 3292
rect 9263 3236 9319 3292
rect 9319 3236 9323 3292
rect 9259 3232 9323 3236
rect 9339 3292 9403 3296
rect 9339 3236 9343 3292
rect 9343 3236 9399 3292
rect 9399 3236 9403 3292
rect 9339 3232 9403 3236
rect 9419 3292 9483 3296
rect 9419 3236 9423 3292
rect 9423 3236 9479 3292
rect 9479 3236 9483 3292
rect 9419 3232 9483 3236
rect 9499 3292 9563 3296
rect 9499 3236 9503 3292
rect 9503 3236 9559 3292
rect 9559 3236 9563 3292
rect 9499 3232 9563 3236
rect 12318 3292 12382 3296
rect 12318 3236 12322 3292
rect 12322 3236 12378 3292
rect 12378 3236 12382 3292
rect 12318 3232 12382 3236
rect 12398 3292 12462 3296
rect 12398 3236 12402 3292
rect 12402 3236 12458 3292
rect 12458 3236 12462 3292
rect 12398 3232 12462 3236
rect 12478 3292 12542 3296
rect 12478 3236 12482 3292
rect 12482 3236 12538 3292
rect 12538 3236 12542 3292
rect 12478 3232 12542 3236
rect 12558 3292 12622 3296
rect 12558 3236 12562 3292
rect 12562 3236 12618 3292
rect 12618 3236 12622 3292
rect 12558 3232 12622 3236
rect 2481 2748 2545 2752
rect 2481 2692 2485 2748
rect 2485 2692 2541 2748
rect 2541 2692 2545 2748
rect 2481 2688 2545 2692
rect 2561 2748 2625 2752
rect 2561 2692 2565 2748
rect 2565 2692 2621 2748
rect 2621 2692 2625 2748
rect 2561 2688 2625 2692
rect 2641 2748 2705 2752
rect 2641 2692 2645 2748
rect 2645 2692 2701 2748
rect 2701 2692 2705 2748
rect 2641 2688 2705 2692
rect 2721 2748 2785 2752
rect 2721 2692 2725 2748
rect 2725 2692 2781 2748
rect 2781 2692 2785 2748
rect 2721 2688 2785 2692
rect 5540 2748 5604 2752
rect 5540 2692 5544 2748
rect 5544 2692 5600 2748
rect 5600 2692 5604 2748
rect 5540 2688 5604 2692
rect 5620 2748 5684 2752
rect 5620 2692 5624 2748
rect 5624 2692 5680 2748
rect 5680 2692 5684 2748
rect 5620 2688 5684 2692
rect 5700 2748 5764 2752
rect 5700 2692 5704 2748
rect 5704 2692 5760 2748
rect 5760 2692 5764 2748
rect 5700 2688 5764 2692
rect 5780 2748 5844 2752
rect 5780 2692 5784 2748
rect 5784 2692 5840 2748
rect 5840 2692 5844 2748
rect 5780 2688 5844 2692
rect 8599 2748 8663 2752
rect 8599 2692 8603 2748
rect 8603 2692 8659 2748
rect 8659 2692 8663 2748
rect 8599 2688 8663 2692
rect 8679 2748 8743 2752
rect 8679 2692 8683 2748
rect 8683 2692 8739 2748
rect 8739 2692 8743 2748
rect 8679 2688 8743 2692
rect 8759 2748 8823 2752
rect 8759 2692 8763 2748
rect 8763 2692 8819 2748
rect 8819 2692 8823 2748
rect 8759 2688 8823 2692
rect 8839 2748 8903 2752
rect 8839 2692 8843 2748
rect 8843 2692 8899 2748
rect 8899 2692 8903 2748
rect 8839 2688 8903 2692
rect 11658 2748 11722 2752
rect 11658 2692 11662 2748
rect 11662 2692 11718 2748
rect 11718 2692 11722 2748
rect 11658 2688 11722 2692
rect 11738 2748 11802 2752
rect 11738 2692 11742 2748
rect 11742 2692 11798 2748
rect 11798 2692 11802 2748
rect 11738 2688 11802 2692
rect 11818 2748 11882 2752
rect 11818 2692 11822 2748
rect 11822 2692 11878 2748
rect 11878 2692 11882 2748
rect 11818 2688 11882 2692
rect 11898 2748 11962 2752
rect 11898 2692 11902 2748
rect 11902 2692 11958 2748
rect 11958 2692 11962 2748
rect 11898 2688 11962 2692
rect 3141 2204 3205 2208
rect 3141 2148 3145 2204
rect 3145 2148 3201 2204
rect 3201 2148 3205 2204
rect 3141 2144 3205 2148
rect 3221 2204 3285 2208
rect 3221 2148 3225 2204
rect 3225 2148 3281 2204
rect 3281 2148 3285 2204
rect 3221 2144 3285 2148
rect 3301 2204 3365 2208
rect 3301 2148 3305 2204
rect 3305 2148 3361 2204
rect 3361 2148 3365 2204
rect 3301 2144 3365 2148
rect 3381 2204 3445 2208
rect 3381 2148 3385 2204
rect 3385 2148 3441 2204
rect 3441 2148 3445 2204
rect 3381 2144 3445 2148
rect 6200 2204 6264 2208
rect 6200 2148 6204 2204
rect 6204 2148 6260 2204
rect 6260 2148 6264 2204
rect 6200 2144 6264 2148
rect 6280 2204 6344 2208
rect 6280 2148 6284 2204
rect 6284 2148 6340 2204
rect 6340 2148 6344 2204
rect 6280 2144 6344 2148
rect 6360 2204 6424 2208
rect 6360 2148 6364 2204
rect 6364 2148 6420 2204
rect 6420 2148 6424 2204
rect 6360 2144 6424 2148
rect 6440 2204 6504 2208
rect 6440 2148 6444 2204
rect 6444 2148 6500 2204
rect 6500 2148 6504 2204
rect 6440 2144 6504 2148
rect 9259 2204 9323 2208
rect 9259 2148 9263 2204
rect 9263 2148 9319 2204
rect 9319 2148 9323 2204
rect 9259 2144 9323 2148
rect 9339 2204 9403 2208
rect 9339 2148 9343 2204
rect 9343 2148 9399 2204
rect 9399 2148 9403 2204
rect 9339 2144 9403 2148
rect 9419 2204 9483 2208
rect 9419 2148 9423 2204
rect 9423 2148 9479 2204
rect 9479 2148 9483 2204
rect 9419 2144 9483 2148
rect 9499 2204 9563 2208
rect 9499 2148 9503 2204
rect 9503 2148 9559 2204
rect 9559 2148 9563 2204
rect 9499 2144 9563 2148
rect 12318 2204 12382 2208
rect 12318 2148 12322 2204
rect 12322 2148 12378 2204
rect 12378 2148 12382 2204
rect 12318 2144 12382 2148
rect 12398 2204 12462 2208
rect 12398 2148 12402 2204
rect 12402 2148 12458 2204
rect 12458 2148 12462 2204
rect 12398 2144 12462 2148
rect 12478 2204 12542 2208
rect 12478 2148 12482 2204
rect 12482 2148 12538 2204
rect 12538 2148 12542 2204
rect 12478 2144 12542 2148
rect 12558 2204 12622 2208
rect 12558 2148 12562 2204
rect 12562 2148 12618 2204
rect 12618 2148 12622 2204
rect 12558 2144 12622 2148
<< metal4 >>
rect 2473 13632 2793 14192
rect 2473 13568 2481 13632
rect 2545 13568 2561 13632
rect 2625 13568 2641 13632
rect 2705 13568 2721 13632
rect 2785 13568 2793 13632
rect 2473 12762 2793 13568
rect 2473 12544 2515 12762
rect 2751 12544 2793 12762
rect 2473 12480 2481 12544
rect 2545 12480 2561 12526
rect 2625 12480 2641 12526
rect 2705 12480 2721 12526
rect 2785 12480 2793 12544
rect 2473 11456 2793 12480
rect 2473 11392 2481 11456
rect 2545 11392 2561 11456
rect 2625 11392 2641 11456
rect 2705 11392 2721 11456
rect 2785 11392 2793 11456
rect 2473 10368 2793 11392
rect 2473 10304 2481 10368
rect 2545 10304 2561 10368
rect 2625 10304 2641 10368
rect 2705 10304 2721 10368
rect 2785 10304 2793 10368
rect 2473 9771 2793 10304
rect 2473 9535 2515 9771
rect 2751 9535 2793 9771
rect 2473 9280 2793 9535
rect 2473 9216 2481 9280
rect 2545 9216 2561 9280
rect 2625 9216 2641 9280
rect 2705 9216 2721 9280
rect 2785 9216 2793 9280
rect 2473 8192 2793 9216
rect 2473 8128 2481 8192
rect 2545 8128 2561 8192
rect 2625 8128 2641 8192
rect 2705 8128 2721 8192
rect 2785 8128 2793 8192
rect 2473 7104 2793 8128
rect 2473 7040 2481 7104
rect 2545 7040 2561 7104
rect 2625 7040 2641 7104
rect 2705 7040 2721 7104
rect 2785 7040 2793 7104
rect 2473 6780 2793 7040
rect 2473 6544 2515 6780
rect 2751 6544 2793 6780
rect 2473 6016 2793 6544
rect 2473 5952 2481 6016
rect 2545 5952 2561 6016
rect 2625 5952 2641 6016
rect 2705 5952 2721 6016
rect 2785 5952 2793 6016
rect 2473 4928 2793 5952
rect 2473 4864 2481 4928
rect 2545 4864 2561 4928
rect 2625 4864 2641 4928
rect 2705 4864 2721 4928
rect 2785 4864 2793 4928
rect 2473 3840 2793 4864
rect 2473 3776 2481 3840
rect 2545 3789 2561 3840
rect 2625 3789 2641 3840
rect 2705 3789 2721 3840
rect 2785 3776 2793 3840
rect 2473 3553 2515 3776
rect 2751 3553 2793 3776
rect 2473 2752 2793 3553
rect 2473 2688 2481 2752
rect 2545 2688 2561 2752
rect 2625 2688 2641 2752
rect 2705 2688 2721 2752
rect 2785 2688 2793 2752
rect 2473 2128 2793 2688
rect 3133 14176 3453 14192
rect 3133 14112 3141 14176
rect 3205 14112 3221 14176
rect 3285 14112 3301 14176
rect 3365 14112 3381 14176
rect 3445 14112 3453 14176
rect 3133 13422 3453 14112
rect 3133 13186 3175 13422
rect 3411 13186 3453 13422
rect 3133 13088 3453 13186
rect 3133 13024 3141 13088
rect 3205 13024 3221 13088
rect 3285 13024 3301 13088
rect 3365 13024 3381 13088
rect 3445 13024 3453 13088
rect 3133 12000 3453 13024
rect 3133 11936 3141 12000
rect 3205 11936 3221 12000
rect 3285 11936 3301 12000
rect 3365 11936 3381 12000
rect 3445 11936 3453 12000
rect 3133 10912 3453 11936
rect 3133 10848 3141 10912
rect 3205 10848 3221 10912
rect 3285 10848 3301 10912
rect 3365 10848 3381 10912
rect 3445 10848 3453 10912
rect 3133 10431 3453 10848
rect 3133 10195 3175 10431
rect 3411 10195 3453 10431
rect 3133 9824 3453 10195
rect 3133 9760 3141 9824
rect 3205 9760 3221 9824
rect 3285 9760 3301 9824
rect 3365 9760 3381 9824
rect 3445 9760 3453 9824
rect 3133 8736 3453 9760
rect 3133 8672 3141 8736
rect 3205 8672 3221 8736
rect 3285 8672 3301 8736
rect 3365 8672 3381 8736
rect 3445 8672 3453 8736
rect 3133 7648 3453 8672
rect 3133 7584 3141 7648
rect 3205 7584 3221 7648
rect 3285 7584 3301 7648
rect 3365 7584 3381 7648
rect 3445 7584 3453 7648
rect 3133 7440 3453 7584
rect 3133 7204 3175 7440
rect 3411 7204 3453 7440
rect 3133 6560 3453 7204
rect 3133 6496 3141 6560
rect 3205 6496 3221 6560
rect 3285 6496 3301 6560
rect 3365 6496 3381 6560
rect 3445 6496 3453 6560
rect 3133 5472 3453 6496
rect 3133 5408 3141 5472
rect 3205 5408 3221 5472
rect 3285 5408 3301 5472
rect 3365 5408 3381 5472
rect 3445 5408 3453 5472
rect 3133 4449 3453 5408
rect 3133 4384 3175 4449
rect 3411 4384 3453 4449
rect 3133 4320 3141 4384
rect 3445 4320 3453 4384
rect 3133 4213 3175 4320
rect 3411 4213 3453 4320
rect 3133 3296 3453 4213
rect 3133 3232 3141 3296
rect 3205 3232 3221 3296
rect 3285 3232 3301 3296
rect 3365 3232 3381 3296
rect 3445 3232 3453 3296
rect 3133 2208 3453 3232
rect 3133 2144 3141 2208
rect 3205 2144 3221 2208
rect 3285 2144 3301 2208
rect 3365 2144 3381 2208
rect 3445 2144 3453 2208
rect 3133 2128 3453 2144
rect 5532 13632 5852 14192
rect 5532 13568 5540 13632
rect 5604 13568 5620 13632
rect 5684 13568 5700 13632
rect 5764 13568 5780 13632
rect 5844 13568 5852 13632
rect 5532 12762 5852 13568
rect 5532 12544 5574 12762
rect 5810 12544 5852 12762
rect 5532 12480 5540 12544
rect 5604 12480 5620 12526
rect 5684 12480 5700 12526
rect 5764 12480 5780 12526
rect 5844 12480 5852 12544
rect 5532 11456 5852 12480
rect 5532 11392 5540 11456
rect 5604 11392 5620 11456
rect 5684 11392 5700 11456
rect 5764 11392 5780 11456
rect 5844 11392 5852 11456
rect 5532 10368 5852 11392
rect 5532 10304 5540 10368
rect 5604 10304 5620 10368
rect 5684 10304 5700 10368
rect 5764 10304 5780 10368
rect 5844 10304 5852 10368
rect 5532 9771 5852 10304
rect 5532 9535 5574 9771
rect 5810 9535 5852 9771
rect 5532 9280 5852 9535
rect 5532 9216 5540 9280
rect 5604 9216 5620 9280
rect 5684 9216 5700 9280
rect 5764 9216 5780 9280
rect 5844 9216 5852 9280
rect 5532 8192 5852 9216
rect 5532 8128 5540 8192
rect 5604 8128 5620 8192
rect 5684 8128 5700 8192
rect 5764 8128 5780 8192
rect 5844 8128 5852 8192
rect 5532 7104 5852 8128
rect 5532 7040 5540 7104
rect 5604 7040 5620 7104
rect 5684 7040 5700 7104
rect 5764 7040 5780 7104
rect 5844 7040 5852 7104
rect 5532 6780 5852 7040
rect 5532 6544 5574 6780
rect 5810 6544 5852 6780
rect 5532 6016 5852 6544
rect 5532 5952 5540 6016
rect 5604 5952 5620 6016
rect 5684 5952 5700 6016
rect 5764 5952 5780 6016
rect 5844 5952 5852 6016
rect 5532 4928 5852 5952
rect 5532 4864 5540 4928
rect 5604 4864 5620 4928
rect 5684 4864 5700 4928
rect 5764 4864 5780 4928
rect 5844 4864 5852 4928
rect 5532 3840 5852 4864
rect 5532 3776 5540 3840
rect 5604 3789 5620 3840
rect 5684 3789 5700 3840
rect 5764 3789 5780 3840
rect 5844 3776 5852 3840
rect 5532 3553 5574 3776
rect 5810 3553 5852 3776
rect 5532 2752 5852 3553
rect 5532 2688 5540 2752
rect 5604 2688 5620 2752
rect 5684 2688 5700 2752
rect 5764 2688 5780 2752
rect 5844 2688 5852 2752
rect 5532 2128 5852 2688
rect 6192 14176 6512 14192
rect 6192 14112 6200 14176
rect 6264 14112 6280 14176
rect 6344 14112 6360 14176
rect 6424 14112 6440 14176
rect 6504 14112 6512 14176
rect 6192 13422 6512 14112
rect 6192 13186 6234 13422
rect 6470 13186 6512 13422
rect 6192 13088 6512 13186
rect 6192 13024 6200 13088
rect 6264 13024 6280 13088
rect 6344 13024 6360 13088
rect 6424 13024 6440 13088
rect 6504 13024 6512 13088
rect 6192 12000 6512 13024
rect 6192 11936 6200 12000
rect 6264 11936 6280 12000
rect 6344 11936 6360 12000
rect 6424 11936 6440 12000
rect 6504 11936 6512 12000
rect 6192 10912 6512 11936
rect 6192 10848 6200 10912
rect 6264 10848 6280 10912
rect 6344 10848 6360 10912
rect 6424 10848 6440 10912
rect 6504 10848 6512 10912
rect 6192 10431 6512 10848
rect 6192 10195 6234 10431
rect 6470 10195 6512 10431
rect 6192 9824 6512 10195
rect 6192 9760 6200 9824
rect 6264 9760 6280 9824
rect 6344 9760 6360 9824
rect 6424 9760 6440 9824
rect 6504 9760 6512 9824
rect 6192 8736 6512 9760
rect 6192 8672 6200 8736
rect 6264 8672 6280 8736
rect 6344 8672 6360 8736
rect 6424 8672 6440 8736
rect 6504 8672 6512 8736
rect 6192 7648 6512 8672
rect 6192 7584 6200 7648
rect 6264 7584 6280 7648
rect 6344 7584 6360 7648
rect 6424 7584 6440 7648
rect 6504 7584 6512 7648
rect 6192 7440 6512 7584
rect 6192 7204 6234 7440
rect 6470 7204 6512 7440
rect 6192 6560 6512 7204
rect 6192 6496 6200 6560
rect 6264 6496 6280 6560
rect 6344 6496 6360 6560
rect 6424 6496 6440 6560
rect 6504 6496 6512 6560
rect 6192 5472 6512 6496
rect 6192 5408 6200 5472
rect 6264 5408 6280 5472
rect 6344 5408 6360 5472
rect 6424 5408 6440 5472
rect 6504 5408 6512 5472
rect 6192 4449 6512 5408
rect 6192 4384 6234 4449
rect 6470 4384 6512 4449
rect 6192 4320 6200 4384
rect 6504 4320 6512 4384
rect 6192 4213 6234 4320
rect 6470 4213 6512 4320
rect 6192 3296 6512 4213
rect 6192 3232 6200 3296
rect 6264 3232 6280 3296
rect 6344 3232 6360 3296
rect 6424 3232 6440 3296
rect 6504 3232 6512 3296
rect 6192 2208 6512 3232
rect 6192 2144 6200 2208
rect 6264 2144 6280 2208
rect 6344 2144 6360 2208
rect 6424 2144 6440 2208
rect 6504 2144 6512 2208
rect 6192 2128 6512 2144
rect 8591 13632 8911 14192
rect 8591 13568 8599 13632
rect 8663 13568 8679 13632
rect 8743 13568 8759 13632
rect 8823 13568 8839 13632
rect 8903 13568 8911 13632
rect 8591 12762 8911 13568
rect 8591 12544 8633 12762
rect 8869 12544 8911 12762
rect 8591 12480 8599 12544
rect 8663 12480 8679 12526
rect 8743 12480 8759 12526
rect 8823 12480 8839 12526
rect 8903 12480 8911 12544
rect 8591 11456 8911 12480
rect 8591 11392 8599 11456
rect 8663 11392 8679 11456
rect 8743 11392 8759 11456
rect 8823 11392 8839 11456
rect 8903 11392 8911 11456
rect 8591 10368 8911 11392
rect 8591 10304 8599 10368
rect 8663 10304 8679 10368
rect 8743 10304 8759 10368
rect 8823 10304 8839 10368
rect 8903 10304 8911 10368
rect 8591 9771 8911 10304
rect 8591 9535 8633 9771
rect 8869 9535 8911 9771
rect 8591 9280 8911 9535
rect 8591 9216 8599 9280
rect 8663 9216 8679 9280
rect 8743 9216 8759 9280
rect 8823 9216 8839 9280
rect 8903 9216 8911 9280
rect 8591 8192 8911 9216
rect 8591 8128 8599 8192
rect 8663 8128 8679 8192
rect 8743 8128 8759 8192
rect 8823 8128 8839 8192
rect 8903 8128 8911 8192
rect 8591 7104 8911 8128
rect 8591 7040 8599 7104
rect 8663 7040 8679 7104
rect 8743 7040 8759 7104
rect 8823 7040 8839 7104
rect 8903 7040 8911 7104
rect 8591 6780 8911 7040
rect 8591 6544 8633 6780
rect 8869 6544 8911 6780
rect 8591 6016 8911 6544
rect 8591 5952 8599 6016
rect 8663 5952 8679 6016
rect 8743 5952 8759 6016
rect 8823 5952 8839 6016
rect 8903 5952 8911 6016
rect 8591 4928 8911 5952
rect 8591 4864 8599 4928
rect 8663 4864 8679 4928
rect 8743 4864 8759 4928
rect 8823 4864 8839 4928
rect 8903 4864 8911 4928
rect 8591 3840 8911 4864
rect 8591 3776 8599 3840
rect 8663 3789 8679 3840
rect 8743 3789 8759 3840
rect 8823 3789 8839 3840
rect 8903 3776 8911 3840
rect 8591 3553 8633 3776
rect 8869 3553 8911 3776
rect 8591 2752 8911 3553
rect 8591 2688 8599 2752
rect 8663 2688 8679 2752
rect 8743 2688 8759 2752
rect 8823 2688 8839 2752
rect 8903 2688 8911 2752
rect 8591 2128 8911 2688
rect 9251 14176 9571 14192
rect 9251 14112 9259 14176
rect 9323 14112 9339 14176
rect 9403 14112 9419 14176
rect 9483 14112 9499 14176
rect 9563 14112 9571 14176
rect 9251 13422 9571 14112
rect 9251 13186 9293 13422
rect 9529 13186 9571 13422
rect 9251 13088 9571 13186
rect 9251 13024 9259 13088
rect 9323 13024 9339 13088
rect 9403 13024 9419 13088
rect 9483 13024 9499 13088
rect 9563 13024 9571 13088
rect 9251 12000 9571 13024
rect 9251 11936 9259 12000
rect 9323 11936 9339 12000
rect 9403 11936 9419 12000
rect 9483 11936 9499 12000
rect 9563 11936 9571 12000
rect 9251 10912 9571 11936
rect 9251 10848 9259 10912
rect 9323 10848 9339 10912
rect 9403 10848 9419 10912
rect 9483 10848 9499 10912
rect 9563 10848 9571 10912
rect 9251 10431 9571 10848
rect 9251 10195 9293 10431
rect 9529 10195 9571 10431
rect 9251 9824 9571 10195
rect 9251 9760 9259 9824
rect 9323 9760 9339 9824
rect 9403 9760 9419 9824
rect 9483 9760 9499 9824
rect 9563 9760 9571 9824
rect 9251 8736 9571 9760
rect 9251 8672 9259 8736
rect 9323 8672 9339 8736
rect 9403 8672 9419 8736
rect 9483 8672 9499 8736
rect 9563 8672 9571 8736
rect 9251 7648 9571 8672
rect 9251 7584 9259 7648
rect 9323 7584 9339 7648
rect 9403 7584 9419 7648
rect 9483 7584 9499 7648
rect 9563 7584 9571 7648
rect 9251 7440 9571 7584
rect 9251 7204 9293 7440
rect 9529 7204 9571 7440
rect 9251 6560 9571 7204
rect 9251 6496 9259 6560
rect 9323 6496 9339 6560
rect 9403 6496 9419 6560
rect 9483 6496 9499 6560
rect 9563 6496 9571 6560
rect 9251 5472 9571 6496
rect 9251 5408 9259 5472
rect 9323 5408 9339 5472
rect 9403 5408 9419 5472
rect 9483 5408 9499 5472
rect 9563 5408 9571 5472
rect 9251 4449 9571 5408
rect 9251 4384 9293 4449
rect 9529 4384 9571 4449
rect 9251 4320 9259 4384
rect 9563 4320 9571 4384
rect 9251 4213 9293 4320
rect 9529 4213 9571 4320
rect 9251 3296 9571 4213
rect 9251 3232 9259 3296
rect 9323 3232 9339 3296
rect 9403 3232 9419 3296
rect 9483 3232 9499 3296
rect 9563 3232 9571 3296
rect 9251 2208 9571 3232
rect 9251 2144 9259 2208
rect 9323 2144 9339 2208
rect 9403 2144 9419 2208
rect 9483 2144 9499 2208
rect 9563 2144 9571 2208
rect 9251 2128 9571 2144
rect 11650 13632 11970 14192
rect 11650 13568 11658 13632
rect 11722 13568 11738 13632
rect 11802 13568 11818 13632
rect 11882 13568 11898 13632
rect 11962 13568 11970 13632
rect 11650 12762 11970 13568
rect 11650 12544 11692 12762
rect 11928 12544 11970 12762
rect 11650 12480 11658 12544
rect 11722 12480 11738 12526
rect 11802 12480 11818 12526
rect 11882 12480 11898 12526
rect 11962 12480 11970 12544
rect 11650 11456 11970 12480
rect 11650 11392 11658 11456
rect 11722 11392 11738 11456
rect 11802 11392 11818 11456
rect 11882 11392 11898 11456
rect 11962 11392 11970 11456
rect 11650 10368 11970 11392
rect 11650 10304 11658 10368
rect 11722 10304 11738 10368
rect 11802 10304 11818 10368
rect 11882 10304 11898 10368
rect 11962 10304 11970 10368
rect 11650 9771 11970 10304
rect 11650 9535 11692 9771
rect 11928 9535 11970 9771
rect 11650 9280 11970 9535
rect 11650 9216 11658 9280
rect 11722 9216 11738 9280
rect 11802 9216 11818 9280
rect 11882 9216 11898 9280
rect 11962 9216 11970 9280
rect 11650 8192 11970 9216
rect 11650 8128 11658 8192
rect 11722 8128 11738 8192
rect 11802 8128 11818 8192
rect 11882 8128 11898 8192
rect 11962 8128 11970 8192
rect 11650 7104 11970 8128
rect 11650 7040 11658 7104
rect 11722 7040 11738 7104
rect 11802 7040 11818 7104
rect 11882 7040 11898 7104
rect 11962 7040 11970 7104
rect 11650 6780 11970 7040
rect 11650 6544 11692 6780
rect 11928 6544 11970 6780
rect 11650 6016 11970 6544
rect 11650 5952 11658 6016
rect 11722 5952 11738 6016
rect 11802 5952 11818 6016
rect 11882 5952 11898 6016
rect 11962 5952 11970 6016
rect 11650 4928 11970 5952
rect 11650 4864 11658 4928
rect 11722 4864 11738 4928
rect 11802 4864 11818 4928
rect 11882 4864 11898 4928
rect 11962 4864 11970 4928
rect 11650 3840 11970 4864
rect 11650 3776 11658 3840
rect 11722 3789 11738 3840
rect 11802 3789 11818 3840
rect 11882 3789 11898 3840
rect 11962 3776 11970 3840
rect 11650 3553 11692 3776
rect 11928 3553 11970 3776
rect 11650 2752 11970 3553
rect 11650 2688 11658 2752
rect 11722 2688 11738 2752
rect 11802 2688 11818 2752
rect 11882 2688 11898 2752
rect 11962 2688 11970 2752
rect 11650 2128 11970 2688
rect 12310 14176 12630 14192
rect 12310 14112 12318 14176
rect 12382 14112 12398 14176
rect 12462 14112 12478 14176
rect 12542 14112 12558 14176
rect 12622 14112 12630 14176
rect 12310 13422 12630 14112
rect 12310 13186 12352 13422
rect 12588 13186 12630 13422
rect 12310 13088 12630 13186
rect 12310 13024 12318 13088
rect 12382 13024 12398 13088
rect 12462 13024 12478 13088
rect 12542 13024 12558 13088
rect 12622 13024 12630 13088
rect 12310 12000 12630 13024
rect 12310 11936 12318 12000
rect 12382 11936 12398 12000
rect 12462 11936 12478 12000
rect 12542 11936 12558 12000
rect 12622 11936 12630 12000
rect 12310 10912 12630 11936
rect 12310 10848 12318 10912
rect 12382 10848 12398 10912
rect 12462 10848 12478 10912
rect 12542 10848 12558 10912
rect 12622 10848 12630 10912
rect 12310 10431 12630 10848
rect 12310 10195 12352 10431
rect 12588 10195 12630 10431
rect 12310 9824 12630 10195
rect 12310 9760 12318 9824
rect 12382 9760 12398 9824
rect 12462 9760 12478 9824
rect 12542 9760 12558 9824
rect 12622 9760 12630 9824
rect 12310 8736 12630 9760
rect 12310 8672 12318 8736
rect 12382 8672 12398 8736
rect 12462 8672 12478 8736
rect 12542 8672 12558 8736
rect 12622 8672 12630 8736
rect 12310 7648 12630 8672
rect 12310 7584 12318 7648
rect 12382 7584 12398 7648
rect 12462 7584 12478 7648
rect 12542 7584 12558 7648
rect 12622 7584 12630 7648
rect 12310 7440 12630 7584
rect 12310 7204 12352 7440
rect 12588 7204 12630 7440
rect 12310 6560 12630 7204
rect 12310 6496 12318 6560
rect 12382 6496 12398 6560
rect 12462 6496 12478 6560
rect 12542 6496 12558 6560
rect 12622 6496 12630 6560
rect 12310 5472 12630 6496
rect 12310 5408 12318 5472
rect 12382 5408 12398 5472
rect 12462 5408 12478 5472
rect 12542 5408 12558 5472
rect 12622 5408 12630 5472
rect 12310 4449 12630 5408
rect 12310 4384 12352 4449
rect 12588 4384 12630 4449
rect 12310 4320 12318 4384
rect 12622 4320 12630 4384
rect 12310 4213 12352 4320
rect 12588 4213 12630 4320
rect 12310 3296 12630 4213
rect 12310 3232 12318 3296
rect 12382 3232 12398 3296
rect 12462 3232 12478 3296
rect 12542 3232 12558 3296
rect 12622 3232 12630 3296
rect 12310 2208 12630 3232
rect 12310 2144 12318 2208
rect 12382 2144 12398 2208
rect 12462 2144 12478 2208
rect 12542 2144 12558 2208
rect 12622 2144 12630 2208
rect 12310 2128 12630 2144
<< via4 >>
rect 2515 12544 2751 12762
rect 2515 12526 2545 12544
rect 2545 12526 2561 12544
rect 2561 12526 2625 12544
rect 2625 12526 2641 12544
rect 2641 12526 2705 12544
rect 2705 12526 2721 12544
rect 2721 12526 2751 12544
rect 2515 9535 2751 9771
rect 2515 6544 2751 6780
rect 2515 3776 2545 3789
rect 2545 3776 2561 3789
rect 2561 3776 2625 3789
rect 2625 3776 2641 3789
rect 2641 3776 2705 3789
rect 2705 3776 2721 3789
rect 2721 3776 2751 3789
rect 2515 3553 2751 3776
rect 3175 13186 3411 13422
rect 3175 10195 3411 10431
rect 3175 7204 3411 7440
rect 3175 4384 3411 4449
rect 3175 4320 3205 4384
rect 3205 4320 3221 4384
rect 3221 4320 3285 4384
rect 3285 4320 3301 4384
rect 3301 4320 3365 4384
rect 3365 4320 3381 4384
rect 3381 4320 3411 4384
rect 3175 4213 3411 4320
rect 5574 12544 5810 12762
rect 5574 12526 5604 12544
rect 5604 12526 5620 12544
rect 5620 12526 5684 12544
rect 5684 12526 5700 12544
rect 5700 12526 5764 12544
rect 5764 12526 5780 12544
rect 5780 12526 5810 12544
rect 5574 9535 5810 9771
rect 5574 6544 5810 6780
rect 5574 3776 5604 3789
rect 5604 3776 5620 3789
rect 5620 3776 5684 3789
rect 5684 3776 5700 3789
rect 5700 3776 5764 3789
rect 5764 3776 5780 3789
rect 5780 3776 5810 3789
rect 5574 3553 5810 3776
rect 6234 13186 6470 13422
rect 6234 10195 6470 10431
rect 6234 7204 6470 7440
rect 6234 4384 6470 4449
rect 6234 4320 6264 4384
rect 6264 4320 6280 4384
rect 6280 4320 6344 4384
rect 6344 4320 6360 4384
rect 6360 4320 6424 4384
rect 6424 4320 6440 4384
rect 6440 4320 6470 4384
rect 6234 4213 6470 4320
rect 8633 12544 8869 12762
rect 8633 12526 8663 12544
rect 8663 12526 8679 12544
rect 8679 12526 8743 12544
rect 8743 12526 8759 12544
rect 8759 12526 8823 12544
rect 8823 12526 8839 12544
rect 8839 12526 8869 12544
rect 8633 9535 8869 9771
rect 8633 6544 8869 6780
rect 8633 3776 8663 3789
rect 8663 3776 8679 3789
rect 8679 3776 8743 3789
rect 8743 3776 8759 3789
rect 8759 3776 8823 3789
rect 8823 3776 8839 3789
rect 8839 3776 8869 3789
rect 8633 3553 8869 3776
rect 9293 13186 9529 13422
rect 9293 10195 9529 10431
rect 9293 7204 9529 7440
rect 9293 4384 9529 4449
rect 9293 4320 9323 4384
rect 9323 4320 9339 4384
rect 9339 4320 9403 4384
rect 9403 4320 9419 4384
rect 9419 4320 9483 4384
rect 9483 4320 9499 4384
rect 9499 4320 9529 4384
rect 9293 4213 9529 4320
rect 11692 12544 11928 12762
rect 11692 12526 11722 12544
rect 11722 12526 11738 12544
rect 11738 12526 11802 12544
rect 11802 12526 11818 12544
rect 11818 12526 11882 12544
rect 11882 12526 11898 12544
rect 11898 12526 11928 12544
rect 11692 9535 11928 9771
rect 11692 6544 11928 6780
rect 11692 3776 11722 3789
rect 11722 3776 11738 3789
rect 11738 3776 11802 3789
rect 11802 3776 11818 3789
rect 11818 3776 11882 3789
rect 11882 3776 11898 3789
rect 11898 3776 11928 3789
rect 11692 3553 11928 3776
rect 12352 13186 12588 13422
rect 12352 10195 12588 10431
rect 12352 7204 12588 7440
rect 12352 4384 12588 4449
rect 12352 4320 12382 4384
rect 12382 4320 12398 4384
rect 12398 4320 12462 4384
rect 12462 4320 12478 4384
rect 12478 4320 12542 4384
rect 12542 4320 12558 4384
rect 12558 4320 12588 4384
rect 12352 4213 12588 4320
<< metal5 >>
rect 1056 13422 13388 13464
rect 1056 13186 3175 13422
rect 3411 13186 6234 13422
rect 6470 13186 9293 13422
rect 9529 13186 12352 13422
rect 12588 13186 13388 13422
rect 1056 13144 13388 13186
rect 1056 12762 13388 12804
rect 1056 12526 2515 12762
rect 2751 12526 5574 12762
rect 5810 12526 8633 12762
rect 8869 12526 11692 12762
rect 11928 12526 13388 12762
rect 1056 12484 13388 12526
rect 1056 10431 13388 10473
rect 1056 10195 3175 10431
rect 3411 10195 6234 10431
rect 6470 10195 9293 10431
rect 9529 10195 12352 10431
rect 12588 10195 13388 10431
rect 1056 10153 13388 10195
rect 1056 9771 13388 9813
rect 1056 9535 2515 9771
rect 2751 9535 5574 9771
rect 5810 9535 8633 9771
rect 8869 9535 11692 9771
rect 11928 9535 13388 9771
rect 1056 9493 13388 9535
rect 1056 7440 13388 7482
rect 1056 7204 3175 7440
rect 3411 7204 6234 7440
rect 6470 7204 9293 7440
rect 9529 7204 12352 7440
rect 12588 7204 13388 7440
rect 1056 7162 13388 7204
rect 1056 6780 13388 6822
rect 1056 6544 2515 6780
rect 2751 6544 5574 6780
rect 5810 6544 8633 6780
rect 8869 6544 11692 6780
rect 11928 6544 13388 6780
rect 1056 6502 13388 6544
rect 1056 4449 13388 4491
rect 1056 4213 3175 4449
rect 3411 4213 6234 4449
rect 6470 4213 9293 4449
rect 9529 4213 12352 4449
rect 12588 4213 13388 4449
rect 1056 4171 13388 4213
rect 1056 3789 13388 3831
rect 1056 3553 2515 3789
rect 2751 3553 5574 3789
rect 5810 3553 8633 3789
rect 8869 3553 11692 3789
rect 11928 3553 13388 3789
rect 1056 3511 13388 3553
use sky130_fd_sc_hd__inv_2  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12144 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1688980957
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1688980957
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1688980957
transform -1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1688980957
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _167_
timestamp 1688980957
transform 1 0 10396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _168_
timestamp 1688980957
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1688980957
transform -1 0 12696 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _172_
timestamp 1688980957
transform -1 0 12052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1688980957
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _176_
timestamp 1688980957
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8556 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7452 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _183_
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _184_
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _185_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _187_
timestamp 1688980957
transform 1 0 6992 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _188_
timestamp 1688980957
transform 1 0 7176 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1688980957
transform -1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1688980957
transform -1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1688980957
transform 1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _194_
timestamp 1688980957
transform 1 0 5888 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _195_
timestamp 1688980957
transform -1 0 6900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _197_
timestamp 1688980957
transform -1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _200_
timestamp 1688980957
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _201_
timestamp 1688980957
transform 1 0 6716 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _203_
timestamp 1688980957
transform -1 0 3496 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _205_
timestamp 1688980957
transform -1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _206_
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _210_
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1688980957
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1688980957
transform -1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _213_
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _214_
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _215_
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _216_
timestamp 1688980957
transform -1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _219_
timestamp 1688980957
transform 1 0 3680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _220_
timestamp 1688980957
transform -1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1688980957
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _223_
timestamp 1688980957
transform -1 0 6164 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1688980957
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1688980957
transform -1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1688980957
transform -1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _229_
timestamp 1688980957
transform 1 0 8188 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9200 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9752 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _233_
timestamp 1688980957
transform -1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _234_
timestamp 1688980957
transform 1 0 9568 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp 1688980957
transform -1 0 11224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 1688980957
transform 1 0 10948 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _239_
timestamp 1688980957
transform -1 0 10212 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _240_
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _241_
timestamp 1688980957
transform 1 0 10212 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1688980957
transform -1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _243_
timestamp 1688980957
transform 1 0 7544 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _244_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _245_
timestamp 1688980957
transform -1 0 9752 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1688980957
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _247_
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _248_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1688980957
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 1688980957
transform -1 0 4324 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _251_
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _252_
timestamp 1688980957
transform 1 0 5336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _254_
timestamp 1688980957
transform 1 0 3312 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _255_
timestamp 1688980957
transform 1 0 4140 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _256_
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1688980957
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _258_
timestamp 1688980957
transform -1 0 4232 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _259_
timestamp 1688980957
transform -1 0 3404 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1688980957
transform 1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _261_
timestamp 1688980957
transform -1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _263_
timestamp 1688980957
transform -1 0 3956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1688980957
transform 1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1688980957
transform -1 0 3036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _267_
timestamp 1688980957
transform -1 0 3312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _268_
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _269_
timestamp 1688980957
transform -1 0 2576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _271_
timestamp 1688980957
transform 1 0 9844 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _272_
timestamp 1688980957
transform 1 0 9108 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10028 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _274_
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _275_
timestamp 1688980957
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _276_
timestamp 1688980957
transform -1 0 4968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _277_
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _278_
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _279_
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _280_
timestamp 1688980957
transform -1 0 5152 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _281_
timestamp 1688980957
transform 1 0 5060 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _282_
timestamp 1688980957
transform 1 0 5888 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _283_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _285_
timestamp 1688980957
transform -1 0 8832 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1688980957
transform -1 0 8004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _287_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _288_
timestamp 1688980957
transform 1 0 8004 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _289_
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _291_
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1688980957
transform -1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1688980957
transform -1 0 3496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1688980957
transform -1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1688980957
transform -1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1688980957
transform -1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1688980957
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1688980957
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1688980957
transform -1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _303_
timestamp 1688980957
transform 1 0 2668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1688980957
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1688980957
transform 1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1688980957
transform 1 0 12144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1688980957
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1688980957
transform 1 0 8464 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1688980957
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1688980957
transform -1 0 8280 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1688980957
transform 1 0 7728 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _319_
timestamp 1688980957
transform 1 0 2576 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _320_
timestamp 1688980957
transform 1 0 1472 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _321_
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1688980957
transform 1 0 5520 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _323_
timestamp 1688980957
transform -1 0 9108 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _328_
timestamp 1688980957
transform 1 0 5060 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _330_
timestamp 1688980957
transform 1 0 5060 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _331_
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _332_
timestamp 1688980957
transform 1 0 10212 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1688980957
transform -1 0 6440 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1688980957
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_48
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_63
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_70
timestamp 1688980957
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_88
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_100
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_123
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_42
timestamp 1688980957
transform 1 0 4968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_64
timestamp 1688980957
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_75
timestamp 1688980957
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_84
timestamp 1688980957
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_94
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_119
timestamp 1688980957
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_126
timestamp 1688980957
transform 1 0 12696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_38
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_59
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_100
timestamp 1688980957
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_104
timestamp 1688980957
transform 1 0 10672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_129
timestamp 1688980957
transform 1 0 12972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_11
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_18
timestamp 1688980957
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_25
timestamp 1688980957
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_34
timestamp 1688980957
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_91
timestamp 1688980957
transform 1 0 9476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_97
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_120
timestamp 1688980957
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_14
timestamp 1688980957
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_23
timestamp 1688980957
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_103
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_107
timestamp 1688980957
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_129
timestamp 1688980957
transform 1 0 12972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_17
timestamp 1688980957
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_25
timestamp 1688980957
transform 1 0 3404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_34
timestamp 1688980957
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1688980957
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_65
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_84
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_90
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_95
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_116
timestamp 1688980957
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_123
timestamp 1688980957
transform 1 0 12420 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_129
timestamp 1688980957
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_11
timestamp 1688980957
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_20
timestamp 1688980957
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_29
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_82
timestamp 1688980957
transform 1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_88
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_101
timestamp 1688980957
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_38
timestamp 1688980957
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_42
timestamp 1688980957
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_68
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_129
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_19
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_31
timestamp 1688980957
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_43
timestamp 1688980957
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_62
timestamp 1688980957
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_87
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 1688980957
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_123
timestamp 1688980957
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_129
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_11
timestamp 1688980957
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_90
timestamp 1688980957
transform 1 0 9384 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_94
timestamp 1688980957
transform 1 0 9752 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_106
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_129
timestamp 1688980957
transform 1 0 12972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_11
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_49
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_77
timestamp 1688980957
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_46
timestamp 1688980957
transform 1 0 5336 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_75
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1688980957
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_114
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_123
timestamp 1688980957
transform 1 0 12420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_129
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_40
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_70
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_101
timestamp 1688980957
transform 1 0 10396 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_120
timestamp 1688980957
transform 1 0 12144 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_21
timestamp 1688980957
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1688980957
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_69
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_107
timestamp 1688980957
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_111
timestamp 1688980957
transform 1 0 11316 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_126
timestamp 1688980957
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_35
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_41
timestamp 1688980957
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_49
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_63
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_89
timestamp 1688980957
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_102
timestamp 1688980957
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_59
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_69
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_75
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_111
timestamp 1688980957
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_123
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_129
timestamp 1688980957
transform 1 0 12972 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_41
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_68
timestamp 1688980957
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_80
timestamp 1688980957
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_102
timestamp 1688980957
transform 1 0 10488 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_123
timestamp 1688980957
transform 1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_129
timestamp 1688980957
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_64
timestamp 1688980957
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_71
timestamp 1688980957
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_119
timestamp 1688980957
transform 1 0 12052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_127
timestamp 1688980957
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_47
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_62
timestamp 1688980957
transform 1 0 6808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_90
timestamp 1688980957
transform 1 0 9384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_97
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_116
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_70
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_90
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_96
timestamp 1688980957
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_120
timestamp 1688980957
transform 1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_128
timestamp 1688980957
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_35
timestamp 1688980957
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1688980957
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_85
timestamp 1688980957
transform 1 0 8924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_97
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 13064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 13064 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform -1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1688980957
transform -1 0 13064 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1688980957
transform -1 0 13064 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1688980957
transform -1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4324 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 3680 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
<< labels >>
flabel metal4 s 3133 2128 3453 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6192 2128 6512 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9251 2128 9571 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12310 2128 12630 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4171 13388 4491 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7162 13388 7482 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10153 13388 10473 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13144 13388 13464 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2473 2128 2793 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5532 2128 5852 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8591 2128 8911 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11650 2128 11970 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3511 13388 3831 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6502 13388 6822 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 9493 13388 9813 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12484 13388 12804 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 pulse_count[0]
port 3 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 pulse_count[1]
port 4 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 pulse_count[2]
port 5 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 pulse_count[3]
port 6 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 pulse_count[4]
port 7 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 pulse_count[5]
port 8 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 pulse_count[6]
port 9 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 pulse_count[7]
port 10 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 pulse_count[8]
port 11 nsew signal input
flabel metal3 s 13657 1912 14457 2032 0 FreeSans 480 0 0 0 pulse_period[0]
port 12 nsew signal input
flabel metal3 s 13657 5992 14457 6112 0 FreeSans 480 0 0 0 pulse_period[1]
port 13 nsew signal input
flabel metal3 s 13657 10072 14457 10192 0 FreeSans 480 0 0 0 pulse_period[2]
port 14 nsew signal input
flabel metal3 s 13657 14152 14457 14272 0 FreeSans 480 0 0 0 pulse_period[3]
port 15 nsew signal input
flabel metal2 s 3606 15801 3662 16601 0 FreeSans 224 90 0 0 pwm_out1
port 16 nsew signal tristate
flabel metal2 s 10782 15801 10838 16601 0 FreeSans 224 90 0 0 pwm_out2
port 17 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 rst
port 18 nsew signal input
rlabel metal1 7222 14144 7222 14144 0 VGND
rlabel metal1 7222 13600 7222 13600 0 VPWR
rlabel metal1 6854 9017 6854 9017 0 _000_
rlabel metal1 7551 5610 7551 5610 0 _001_
rlabel metal1 8418 9146 8418 9146 0 _002_
rlabel metal1 3135 6698 3135 6698 0 _003_
rlabel metal1 2583 8874 2583 8874 0 _004_
rlabel metal1 4377 9622 4377 9622 0 _005_
rlabel metal2 2898 5882 2898 5882 0 _006_
rlabel metal1 5842 5338 5842 5338 0 _007_
rlabel metal1 6808 7174 6808 7174 0 _008_
rlabel metal2 8050 7582 8050 7582 0 _009_
rlabel metal1 10902 7310 10902 7310 0 _010_
rlabel metal2 12466 6936 12466 6936 0 _011_
rlabel metal2 12190 4760 12190 4760 0 _012_
rlabel metal1 12650 3162 12650 3162 0 _013_
rlabel metal1 6026 9656 6026 9656 0 _014_
rlabel metal2 4738 10914 4738 10914 0 _015_
rlabel metal1 5842 12750 5842 12750 0 _016_
rlabel metal1 8556 12410 8556 12410 0 _017_
rlabel metal2 11638 13124 11638 13124 0 _018_
rlabel metal1 12466 8296 12466 8296 0 _019_
rlabel metal2 5750 8738 5750 8738 0 _020_
rlabel metal2 8786 5576 8786 5576 0 _021_
rlabel metal1 8234 9486 8234 9486 0 _022_
rlabel metal1 1971 6970 1971 6970 0 _023_
rlabel metal1 3128 8602 3128 8602 0 _024_
rlabel metal1 2944 9622 2944 9622 0 _025_
rlabel metal1 1978 5746 1978 5746 0 _026_
rlabel metal1 4692 6358 4692 6358 0 _027_
rlabel metal1 5927 6970 5927 6970 0 _028_
rlabel metal1 8602 7446 8602 7446 0 _029_
rlabel metal1 9568 7446 9568 7446 0 _030_
rlabel metal1 11270 6698 11270 6698 0 _031_
rlabel metal1 11500 4658 11500 4658 0 _032_
rlabel metal1 12236 3162 12236 3162 0 _033_
rlabel metal1 5658 10098 5658 10098 0 _034_
rlabel metal1 4232 11050 4232 11050 0 _035_
rlabel metal1 5980 12614 5980 12614 0 _036_
rlabel metal1 7820 12750 7820 12750 0 _037_
rlabel metal1 10534 13192 10534 13192 0 _038_
rlabel metal2 11454 8364 11454 8364 0 _039_
rlabel metal1 7176 12886 7176 12886 0 _040_
rlabel metal1 7774 12410 7774 12410 0 _041_
rlabel metal1 8786 13158 8786 13158 0 _042_
rlabel metal1 9522 13294 9522 13294 0 _043_
rlabel via1 7414 12138 7414 12138 0 _044_
rlabel metal1 7590 12308 7590 12308 0 _045_
rlabel metal1 6900 12614 6900 12614 0 _046_
rlabel metal1 6616 12886 6616 12886 0 _047_
rlabel metal1 6256 12818 6256 12818 0 _048_
rlabel metal1 6762 10710 6762 10710 0 _049_
rlabel metal1 6164 10778 6164 10778 0 _050_
rlabel metal1 7314 10778 7314 10778 0 _051_
rlabel metal2 6946 3298 6946 3298 0 _052_
rlabel metal1 7268 3706 7268 3706 0 _053_
rlabel metal1 10425 4114 10425 4114 0 _054_
rlabel metal1 5934 8432 5934 8432 0 _055_
rlabel metal1 2346 8398 2346 8398 0 _056_
rlabel metal1 4692 5270 4692 5270 0 _057_
rlabel metal1 9928 6630 9928 6630 0 _058_
rlabel metal2 9890 6562 9890 6562 0 _059_
rlabel metal1 10994 5236 10994 5236 0 _060_
rlabel metal1 12144 3026 12144 3026 0 _061_
rlabel metal1 11040 4998 11040 4998 0 _062_
rlabel metal1 9890 3502 9890 3502 0 _063_
rlabel metal1 5152 3570 5152 3570 0 _064_
rlabel metal1 4186 3638 4186 3638 0 _065_
rlabel metal1 2944 3162 2944 3162 0 _066_
rlabel metal1 1886 3400 1886 3400 0 _067_
rlabel metal2 3082 3332 3082 3332 0 _068_
rlabel metal1 5014 3434 5014 3434 0 _069_
rlabel metal1 4094 3604 4094 3604 0 _070_
rlabel metal1 4278 3094 4278 3094 0 _071_
rlabel metal1 4370 3060 4370 3060 0 _072_
rlabel metal1 4416 2822 4416 2822 0 _073_
rlabel metal1 6118 3536 6118 3536 0 _074_
rlabel metal1 5382 2958 5382 2958 0 _075_
rlabel metal1 6210 3706 6210 3706 0 _076_
rlabel metal1 7728 3366 7728 3366 0 _077_
rlabel metal1 8878 4046 8878 4046 0 _078_
rlabel metal1 8924 3502 8924 3502 0 _079_
rlabel metal1 8372 3434 8372 3434 0 _080_
rlabel metal1 8970 3162 8970 3162 0 _081_
rlabel metal2 8970 3672 8970 3672 0 _082_
rlabel metal2 9706 3332 9706 3332 0 _083_
rlabel metal1 10948 3706 10948 3706 0 _084_
rlabel metal1 10097 3570 10097 3570 0 _085_
rlabel metal1 10488 3706 10488 3706 0 _086_
rlabel metal1 10810 4012 10810 4012 0 _087_
rlabel metal1 2254 7990 2254 7990 0 _088_
rlabel metal1 11546 5202 11546 5202 0 _089_
rlabel metal1 9752 6630 9752 6630 0 _090_
rlabel metal1 10488 6426 10488 6426 0 _091_
rlabel metal1 10856 6766 10856 6766 0 _092_
rlabel metal1 8510 6766 8510 6766 0 _093_
rlabel metal1 9338 6732 9338 6732 0 _094_
rlabel metal1 9154 6868 9154 6868 0 _095_
rlabel metal1 8510 6426 8510 6426 0 _096_
rlabel metal1 8556 6970 8556 6970 0 _097_
rlabel metal1 4186 6426 4186 6426 0 _098_
rlabel metal1 5704 6698 5704 6698 0 _099_
rlabel metal1 6210 7446 6210 7446 0 _100_
rlabel metal2 3726 5712 3726 5712 0 _101_
rlabel metal1 4462 5610 4462 5610 0 _102_
rlabel metal1 4738 5542 4738 5542 0 _103_
rlabel metal1 3404 5270 3404 5270 0 _104_
rlabel metal1 2691 6290 2691 6290 0 _105_
rlabel metal1 2668 7378 2668 7378 0 _106_
rlabel metal1 3772 8534 3772 8534 0 _107_
rlabel metal1 3496 8602 3496 8602 0 _108_
rlabel metal1 2576 7854 2576 7854 0 _109_
rlabel metal1 2622 8500 2622 8500 0 _110_
rlabel metal1 2576 7514 2576 7514 0 _111_
rlabel metal2 9062 11730 9062 11730 0 _112_
rlabel metal1 9660 11526 9660 11526 0 _113_
rlabel metal2 9706 12614 9706 12614 0 _114_
rlabel metal1 10258 12138 10258 12138 0 _115_
rlabel metal1 9706 10710 9706 10710 0 _116_
rlabel metal1 4692 3162 4692 3162 0 _117_
rlabel metal1 3266 3536 3266 3536 0 _118_
rlabel metal1 3818 3536 3818 3536 0 _119_
rlabel metal1 4692 3706 4692 3706 0 _120_
rlabel metal1 5428 4114 5428 4114 0 _121_
rlabel metal1 5796 3162 5796 3162 0 _122_
rlabel metal1 6026 3638 6026 3638 0 _123_
rlabel metal1 7130 3094 7130 3094 0 _124_
rlabel metal2 7498 3196 7498 3196 0 _125_
rlabel metal1 7774 3060 7774 3060 0 _126_
rlabel metal1 8050 3162 8050 3162 0 _127_
rlabel metal1 8510 3706 8510 3706 0 _128_
rlabel metal1 8556 3910 8556 3910 0 _129_
rlabel metal1 9982 4794 9982 4794 0 _130_
rlabel metal1 3036 6290 3036 6290 0 _131_
rlabel metal1 5658 12784 5658 12784 0 _132_
rlabel metal1 12236 9146 12236 9146 0 _133_
rlabel metal1 7176 10030 7176 10030 0 _134_
rlabel metal1 9246 11152 9246 11152 0 _135_
rlabel metal1 9522 11084 9522 11084 0 _136_
rlabel metal1 10120 12682 10120 12682 0 _137_
rlabel metal2 11178 11424 11178 11424 0 _138_
rlabel metal1 7268 8466 7268 8466 0 _139_
rlabel metal2 9798 10438 9798 10438 0 _140_
rlabel metal1 10166 9894 10166 9894 0 _141_
rlabel metal1 10764 10234 10764 10234 0 _142_
rlabel metal1 11454 10506 11454 10506 0 _143_
rlabel metal1 12098 10098 12098 10098 0 _144_
rlabel metal1 11960 10778 11960 10778 0 _145_
rlabel metal1 12098 10540 12098 10540 0 _146_
rlabel metal1 11454 11662 11454 11662 0 _147_
rlabel metal1 9982 10676 9982 10676 0 _148_
rlabel metal1 12006 11152 12006 11152 0 _149_
rlabel metal1 10764 9622 10764 9622 0 _150_
rlabel metal1 11362 10030 11362 10030 0 _151_
rlabel metal1 12144 10234 12144 10234 0 _152_
rlabel metal1 10074 10608 10074 10608 0 _153_
rlabel metal1 9016 10710 9016 10710 0 _154_
rlabel metal1 6762 12818 6762 12818 0 _155_
rlabel metal1 6394 10642 6394 10642 0 _156_
rlabel metal2 4094 11815 4094 11815 0 clk
rlabel metal1 7360 7854 7360 7854 0 clknet_0_clk
rlabel metal1 1472 5746 1472 5746 0 clknet_1_0__leaf_clk
rlabel metal1 2622 9418 2622 9418 0 clknet_1_1__leaf_clk
rlabel metal1 2346 3638 2346 3638 0 counter1\[0\]
rlabel metal1 12926 4148 12926 4148 0 counter1\[10\]
rlabel metal1 2208 3366 2208 3366 0 counter1\[1\]
rlabel metal1 4311 9010 4311 9010 0 counter1\[2\]
rlabel metal1 4600 4114 4600 4114 0 counter1\[3\]
rlabel metal2 4278 6528 4278 6528 0 counter1\[4\]
rlabel metal2 5566 5389 5566 5389 0 counter1\[5\]
rlabel metal1 7452 6766 7452 6766 0 counter1\[6\]
rlabel metal2 10166 6936 10166 6936 0 counter1\[7\]
rlabel metal1 10304 6358 10304 6358 0 counter1\[8\]
rlabel metal1 11178 4250 11178 4250 0 counter1\[9\]
rlabel metal2 7406 9860 7406 9860 0 counter2\[0\]
rlabel metal1 7222 11084 7222 11084 0 counter2\[1\]
rlabel metal1 9430 12104 9430 12104 0 counter2\[2\]
rlabel metal1 9384 12750 9384 12750 0 counter2\[3\]
rlabel metal1 8418 12240 8418 12240 0 counter2\[4\]
rlabel metal2 12926 8228 12926 8228 0 counter2\[5\]
rlabel metal1 2484 4046 2484 4046 0 net1
rlabel metal1 12972 2618 12972 2618 0 net10
rlabel metal1 11914 9554 11914 9554 0 net11
rlabel metal1 12098 9486 12098 9486 0 net12
rlabel metal1 12420 13770 12420 13770 0 net13
rlabel metal1 2714 4522 2714 4522 0 net14
rlabel metal1 5842 5882 5842 5882 0 net15
rlabel metal2 10994 13163 10994 13163 0 net16
rlabel metal1 6716 8602 6716 8602 0 net17
rlabel metal1 12282 8534 12282 8534 0 net18
rlabel metal1 8096 5134 8096 5134 0 net19
rlabel metal1 2852 2618 2852 2618 0 net2
rlabel metal1 12052 4114 12052 4114 0 net20
rlabel metal1 7912 10642 7912 10642 0 net21
rlabel metal1 4784 2618 4784 2618 0 net3
rlabel metal1 5934 3502 5934 3502 0 net4
rlabel metal1 6486 2584 6486 2584 0 net5
rlabel metal1 8786 3026 8786 3026 0 net6
rlabel metal2 10442 2788 10442 2788 0 net7
rlabel metal1 11454 2482 11454 2482 0 net8
rlabel metal1 12834 2924 12834 2924 0 net9
rlabel metal1 7222 8840 7222 8840 0 prev_pwm_out2
rlabel metal2 966 1588 966 1588 0 pulse_count[0]
rlabel metal2 2530 1588 2530 1588 0 pulse_count[1]
rlabel metal2 4094 1588 4094 1588 0 pulse_count[2]
rlabel metal2 5658 1588 5658 1588 0 pulse_count[3]
rlabel metal2 7222 1588 7222 1588 0 pulse_count[4]
rlabel metal2 8786 1588 8786 1588 0 pulse_count[5]
rlabel metal2 10350 1588 10350 1588 0 pulse_count[6]
rlabel metal2 11914 1554 11914 1554 0 pulse_count[7]
rlabel metal2 13478 1894 13478 1894 0 pulse_count[8]
rlabel metal1 13110 2346 13110 2346 0 pulse_period[0]
rlabel metal2 13018 6137 13018 6137 0 pulse_period[1]
rlabel metal2 13018 10353 13018 10353 0 pulse_period[2]
rlabel metal1 13110 13974 13110 13974 0 pulse_period[3]
rlabel metal1 3772 14042 3772 14042 0 pwm_out1
rlabel metal1 10948 14042 10948 14042 0 pwm_out2
rlabel metal3 820 4148 820 4148 0 rst
<< properties >>
string FIXED_BBOX 0 0 14457 16601
<< end >>
