magic
tech sky130A
magscale 1 2
timestamp 1717264603
<< nwell >>
rect 22439 1246 22473 1301
rect 26848 1245 26882 1279
rect 27024 1245 27058 1279
rect 31268 1245 31302 1302
rect 31444 1245 31478 1302
rect 31220 1166 31221 1182
rect 31020 979 31221 1166
<< poly >>
rect 21005 9050 21035 9060
rect 21005 8794 21035 8813
rect 20646 8764 21035 8794
rect 20646 8758 20753 8764
rect 20646 8671 20656 8758
rect 20743 8671 20753 8758
rect 21343 8726 21373 8808
rect 21431 8772 21765 8803
rect 21343 8696 21493 8726
rect 20646 8655 20753 8671
rect 21463 8667 21493 8696
rect 21544 8669 21610 8679
rect 21734 8676 21765 8772
rect 21544 8667 21560 8669
rect 21463 8637 21560 8667
rect 21544 8635 21560 8637
rect 21594 8635 21610 8669
rect 21544 8625 21610 8635
rect 21723 8660 21777 8676
rect 21723 8626 21733 8660
rect 21767 8626 21777 8660
rect 21723 8610 21777 8626
rect 25040 7542 25118 7565
rect 25040 7508 25062 7542
rect 25096 7508 25118 7542
rect 25040 7486 25118 7508
rect 25508 7439 25558 7495
rect 25506 7423 25560 7439
rect 25506 7389 25516 7423
rect 25550 7389 25560 7423
rect 25506 7373 25560 7389
rect 26859 1526 26913 1542
rect 26859 1492 26869 1526
rect 26903 1492 26913 1526
rect 26859 1476 26913 1492
rect 31263 1522 31317 1538
rect 31263 1488 31273 1522
rect 31307 1488 31317 1522
rect 22457 1456 22523 1472
rect 22457 1422 22473 1456
rect 22507 1422 22523 1456
rect 22457 1406 22523 1422
rect 26871 1417 26901 1476
rect 31263 1472 31317 1488
rect 22475 1364 22505 1406
rect 26758 1387 27012 1417
rect 31275 1405 31305 1472
rect 22374 1334 22603 1364
rect 22374 611 22404 1334
rect 22573 1267 22603 1334
rect 22485 611 22515 626
rect 22374 581 22515 611
rect 22573 594 22603 635
rect 26758 610 26788 1387
rect 26982 1265 27012 1387
rect 31160 1375 31432 1405
rect 26894 610 26924 625
rect 22573 584 22677 594
rect 18124 422 18154 577
rect 22573 552 22627 584
rect 22611 550 22627 552
rect 22661 550 22677 584
rect 26758 580 26924 610
rect 26982 584 27012 625
rect 31160 606 31190 1375
rect 31402 1267 31432 1375
rect 31314 606 31344 634
rect 22611 540 22677 550
rect 26982 574 27086 584
rect 31160 576 31344 606
rect 31402 584 31432 625
rect 26982 542 27036 574
rect 27020 540 27036 542
rect 27070 540 27086 574
rect 31402 574 31506 584
rect 31402 542 31456 574
rect 27020 530 27086 540
rect 31440 540 31456 542
rect 31490 540 31506 574
rect 31440 530 31506 540
rect 18112 406 18166 422
rect 18112 372 18122 406
rect 18156 372 18166 406
rect 18112 356 18166 372
<< polycont >>
rect 20656 8671 20743 8758
rect 21560 8635 21594 8669
rect 21733 8626 21767 8660
rect 25062 7508 25096 7542
rect 25516 7389 25550 7423
rect 26869 1492 26903 1526
rect 31273 1488 31307 1522
rect 22473 1422 22507 1456
rect 22627 550 22661 584
rect 27036 540 27070 574
rect 31456 540 31490 574
rect 18122 372 18156 406
<< locali >>
rect 21087 9496 21121 11197
rect 20640 8671 20646 8758
rect 20753 8671 20759 8758
rect 21560 8669 21594 8685
rect 21560 8619 21594 8635
rect 21717 8626 21733 8660
rect 21767 8626 21783 8660
rect 25040 7550 25118 7565
rect 25040 7500 25054 7550
rect 25104 7500 25118 7550
rect 25040 7486 25118 7500
rect 25500 7389 25508 7423
rect 25558 7389 25566 7423
rect 27083 6025 27239 8328
rect 27071 6012 27252 6025
rect 27071 5856 27083 6012
rect 27239 5856 27252 6012
rect 27071 5843 27252 5856
rect 22374 2003 22408 2004
rect 22374 1301 22408 1969
rect 22457 1422 22473 1456
rect 22507 1422 22523 1456
rect 22374 1267 22473 1301
rect 22439 1246 22473 1267
rect 22615 1246 22649 1967
rect 26755 1331 26789 1950
rect 26853 1492 26869 1526
rect 26903 1492 26919 1526
rect 26755 1297 26882 1331
rect 17462 938 17468 1137
rect 17667 938 18092 1137
rect 26848 1242 26882 1297
rect 27024 1245 27058 1952
rect 31158 1339 31192 2019
rect 31257 1488 31273 1522
rect 31307 1488 31323 1522
rect 31158 1305 31302 1339
rect 22727 1147 22828 1155
rect 27135 1150 27235 1164
rect 31268 1245 31302 1305
rect 31444 1245 31478 1733
rect 30864 1118 30964 1149
rect 16955 794 18081 800
rect 16955 607 16961 794
rect 17148 607 18081 794
rect 22903 829 22989 838
rect 27311 827 27397 881
rect 31040 790 31127 803
rect 18459 732 18545 784
rect 16955 601 18081 607
rect 18086 406 18194 440
rect 18086 372 18122 406
rect 18156 372 18194 406
rect 18086 336 18194 372
rect 22527 340 22561 648
rect 22627 596 22661 600
rect 22615 584 22673 596
rect 22615 550 22627 584
rect 22661 550 22673 584
rect 22615 538 22673 550
rect 22627 534 22661 538
rect 22492 307 22594 340
rect 26936 339 26970 647
rect 27036 586 27070 590
rect 27024 574 27082 586
rect 27024 540 27036 574
rect 27070 540 27082 574
rect 27024 528 27082 540
rect 27036 524 27070 528
rect 31356 339 31390 647
rect 31456 586 31490 590
rect 31444 574 31502 586
rect 31444 540 31456 574
rect 31490 540 31502 574
rect 31444 528 31502 540
rect 31456 524 31490 528
rect 22492 273 22527 307
rect 22561 273 22594 307
rect 22492 244 22594 273
rect 26901 306 27003 339
rect 26901 272 26936 306
rect 26970 272 27003 306
rect 26901 243 27003 272
rect 31321 306 31423 339
rect 31321 272 31356 306
rect 31390 272 31423 306
rect 31321 243 31423 272
<< viali >>
rect 21087 11197 21121 11231
rect 20646 8758 20753 8768
rect 20646 8671 20656 8758
rect 20656 8671 20743 8758
rect 20743 8671 20753 8758
rect 20646 8661 20753 8671
rect 21560 8635 21594 8669
rect 21733 8626 21767 8660
rect 25054 7542 25104 7550
rect 25054 7508 25062 7542
rect 25062 7508 25096 7542
rect 25096 7508 25104 7542
rect 25054 7500 25104 7508
rect 25508 7423 25558 7431
rect 25508 7389 25516 7423
rect 25516 7389 25550 7423
rect 25550 7389 25558 7423
rect 25508 7381 25558 7389
rect 27083 5856 27239 6012
rect 31158 2019 31192 2053
rect 22374 1969 22408 2003
rect 22615 1967 22649 2001
rect 22473 1422 22507 1456
rect 26755 1950 26789 1984
rect 27024 1952 27058 1986
rect 26869 1492 26903 1526
rect 17468 938 17667 1137
rect 18283 1077 18383 1177
rect 22727 1155 22828 1256
rect 31374 1733 31518 1877
rect 31273 1488 31307 1522
rect 27135 1164 27235 1264
rect 30864 1149 30964 1249
rect 16961 607 17148 794
rect 18459 784 18545 870
rect 22903 838 22989 924
rect 27311 881 27397 967
rect 31040 803 31127 890
rect 18122 372 18156 406
rect 22627 550 22661 584
rect 27036 540 27070 574
rect 31456 540 31490 574
rect 22527 273 22561 307
rect 26936 272 26970 306
rect 31356 272 31390 306
<< metal1 >>
rect 19705 30937 20105 33423
rect 19961 11345 20278 11355
rect 19961 11048 19972 11345
rect 20269 11231 24223 11345
rect 20269 11197 21087 11231
rect 21121 11197 24223 11231
rect 20269 11048 24223 11197
rect 19961 11038 20278 11048
rect 20634 8774 20765 8780
rect 20634 8655 20640 8774
rect 20759 8655 20765 8774
rect 20634 8649 20765 8655
rect 21544 8678 21611 8686
rect 21544 8626 21551 8678
rect 21603 8626 21611 8678
rect 21544 8620 21611 8626
rect 21717 8669 21784 8676
rect 21717 8617 21724 8669
rect 21776 8617 21784 8669
rect 21717 8610 21784 8617
rect 19962 6530 20279 6542
rect 21103 6530 21137 8474
rect 25040 7556 25118 7565
rect 25040 7494 25048 7556
rect 25110 7494 25118 7556
rect 25040 7486 25118 7494
rect 25493 7437 25574 7447
rect 25493 7375 25502 7437
rect 25564 7375 25574 7437
rect 25493 7369 25574 7375
rect 19962 6233 19972 6530
rect 20269 6233 24839 6530
rect 19962 6223 20279 6233
rect 27071 6018 27252 6025
rect 27071 5850 27077 6018
rect 27245 5850 27252 6018
rect 27071 5843 27252 5850
rect 25051 5202 25103 5208
rect 22600 5150 22606 5202
rect 22658 5193 22664 5202
rect 22658 5159 25051 5193
rect 22658 5150 22664 5159
rect 25051 5144 25103 5150
rect 22888 4870 22944 4876
rect 26740 4859 26746 4868
rect 22944 4825 26746 4859
rect 26740 4816 26746 4825
rect 26798 4816 26804 4868
rect 22888 4808 22944 4814
rect 23465 4374 23517 4380
rect 31149 4374 31201 4380
rect 23517 4331 31149 4365
rect 23465 4316 23517 4322
rect 31149 4316 31201 4322
rect 31152 2062 31198 2065
rect 22359 2012 22423 2018
rect 22359 1960 22365 2012
rect 22417 1960 22423 2012
rect 22359 1954 22423 1960
rect 22600 2010 22664 2016
rect 31143 2010 31149 2062
rect 31201 2010 31207 2062
rect 22600 1958 22606 2010
rect 22658 1958 22664 2010
rect 31152 2007 31198 2010
rect 22600 1952 22664 1958
rect 26740 1993 26804 1999
rect 26740 1941 26746 1993
rect 26798 1941 26804 1993
rect 26740 1935 26804 1941
rect 27009 1995 27073 2001
rect 27009 1943 27015 1995
rect 27067 1943 27073 1995
rect 27009 1937 27073 1943
rect 31362 1727 31368 1883
rect 31524 1727 31530 1883
rect 18160 1649 31307 1695
rect 17453 1143 17686 1153
rect 17453 932 17462 1143
rect 17673 932 17686 1143
rect 18160 1136 18206 1649
rect 22473 1472 22507 1649
rect 26869 1542 26903 1649
rect 26853 1526 26919 1542
rect 31273 1538 31307 1649
rect 26853 1492 26869 1526
rect 26903 1492 26919 1526
rect 26853 1476 26919 1492
rect 31257 1522 31323 1538
rect 31257 1488 31273 1522
rect 31307 1488 31323 1522
rect 31257 1472 31323 1488
rect 22457 1456 22523 1472
rect 22457 1422 22473 1456
rect 22507 1422 22523 1456
rect 22457 1406 22523 1422
rect 22712 1262 22843 1272
rect 18271 1183 18396 1192
rect 18271 1071 18277 1183
rect 18389 1071 18396 1183
rect 22712 1149 22721 1262
rect 22834 1149 22843 1262
rect 27120 1270 27250 1279
rect 27120 1158 27129 1270
rect 27241 1158 27250 1270
rect 27120 1149 27250 1158
rect 30849 1255 30979 1264
rect 22712 1140 22843 1149
rect 30849 1143 30858 1255
rect 30970 1143 30979 1255
rect 30849 1134 30979 1143
rect 18271 1065 18396 1071
rect 27294 973 27414 984
rect 17453 923 17686 932
rect 22888 930 23004 941
rect 18444 876 18560 887
rect 16949 800 17161 807
rect 16949 601 16955 800
rect 17154 601 17161 800
rect 18444 778 18453 876
rect 18551 778 18560 876
rect 22888 832 22897 930
rect 22995 832 23004 930
rect 27294 875 27305 973
rect 27403 875 27414 973
rect 27294 864 27414 875
rect 31022 896 31144 907
rect 22888 823 23004 832
rect 31022 797 31034 896
rect 31133 797 31144 896
rect 31022 786 31144 797
rect 18444 768 18560 778
rect 16949 595 17161 601
rect 22615 584 22673 596
rect 22615 550 22627 584
rect 22661 550 22673 584
rect 22615 515 22673 550
rect 27024 574 27082 586
rect 27024 540 27036 574
rect 27070 540 27082 574
rect 27024 515 27082 540
rect 31444 574 31502 586
rect 31444 540 31456 574
rect 31490 540 31502 574
rect 31444 515 31502 540
rect 18086 457 31502 515
rect 18086 415 18194 457
rect 18086 363 18113 415
rect 18165 363 18194 415
rect 18086 336 18194 363
rect 22492 316 22594 340
rect 22492 264 22518 316
rect 22570 264 22594 316
rect 22492 244 22594 264
rect 26901 315 27003 339
rect 26901 263 26927 315
rect 26979 263 27003 315
rect 26901 243 27003 263
rect 31321 315 31423 339
rect 31321 263 31347 315
rect 31399 263 31423 315
rect 31321 243 31423 263
<< via1 >>
rect 19972 11048 20269 11345
rect 20640 8768 20759 8774
rect 20640 8661 20646 8768
rect 20646 8661 20753 8768
rect 20753 8661 20759 8768
rect 20640 8655 20759 8661
rect 21551 8669 21603 8678
rect 21551 8635 21560 8669
rect 21560 8635 21594 8669
rect 21594 8635 21603 8669
rect 21551 8626 21603 8635
rect 21724 8660 21776 8669
rect 21724 8626 21733 8660
rect 21733 8626 21767 8660
rect 21767 8626 21776 8660
rect 21724 8617 21776 8626
rect 25048 7550 25110 7556
rect 25048 7500 25054 7550
rect 25054 7500 25104 7550
rect 25104 7500 25110 7550
rect 25048 7494 25110 7500
rect 25502 7431 25564 7437
rect 25502 7381 25508 7431
rect 25508 7381 25558 7431
rect 25558 7381 25564 7431
rect 25502 7375 25564 7381
rect 19972 6233 20269 6530
rect 27077 6012 27245 6018
rect 27077 5856 27083 6012
rect 27083 5856 27239 6012
rect 27239 5856 27245 6012
rect 27077 5850 27245 5856
rect 22606 5150 22658 5202
rect 25051 5150 25103 5202
rect 22888 4814 22944 4870
rect 26746 4816 26798 4868
rect 23465 4322 23517 4374
rect 31149 4322 31201 4374
rect 22365 2003 22417 2012
rect 22365 1969 22374 2003
rect 22374 1969 22408 2003
rect 22408 1969 22417 2003
rect 22365 1960 22417 1969
rect 31149 2053 31201 2062
rect 31149 2019 31158 2053
rect 31158 2019 31192 2053
rect 31192 2019 31201 2053
rect 31149 2010 31201 2019
rect 22606 2001 22658 2010
rect 22606 1967 22615 2001
rect 22615 1967 22649 2001
rect 22649 1967 22658 2001
rect 22606 1958 22658 1967
rect 26746 1984 26798 1993
rect 26746 1950 26755 1984
rect 26755 1950 26789 1984
rect 26789 1950 26798 1984
rect 26746 1941 26798 1950
rect 27015 1986 27067 1995
rect 27015 1952 27024 1986
rect 27024 1952 27058 1986
rect 27058 1952 27067 1986
rect 27015 1943 27067 1952
rect 31368 1877 31524 1883
rect 31368 1733 31374 1877
rect 31374 1733 31518 1877
rect 31518 1733 31524 1877
rect 31368 1727 31524 1733
rect 17462 1137 17673 1143
rect 17462 938 17468 1137
rect 17468 938 17667 1137
rect 17667 938 17673 1137
rect 17462 932 17673 938
rect 18277 1177 18389 1183
rect 18277 1077 18283 1177
rect 18283 1077 18383 1177
rect 18383 1077 18389 1177
rect 18277 1071 18389 1077
rect 22721 1256 22834 1262
rect 22721 1155 22727 1256
rect 22727 1155 22828 1256
rect 22828 1155 22834 1256
rect 22721 1149 22834 1155
rect 27129 1264 27241 1270
rect 27129 1164 27135 1264
rect 27135 1164 27235 1264
rect 27235 1164 27241 1264
rect 27129 1158 27241 1164
rect 30858 1249 30970 1255
rect 30858 1149 30864 1249
rect 30864 1149 30964 1249
rect 30964 1149 30970 1249
rect 30858 1143 30970 1149
rect 16955 794 17154 800
rect 16955 607 16961 794
rect 16961 607 17148 794
rect 17148 607 17154 794
rect 16955 601 17154 607
rect 18453 870 18551 876
rect 18453 784 18459 870
rect 18459 784 18545 870
rect 18545 784 18551 870
rect 18453 778 18551 784
rect 22897 924 22995 930
rect 22897 838 22903 924
rect 22903 838 22989 924
rect 22989 838 22995 924
rect 22897 832 22995 838
rect 27305 967 27403 973
rect 27305 881 27311 967
rect 27311 881 27397 967
rect 27397 881 27403 967
rect 27305 875 27403 881
rect 31034 890 31133 896
rect 31034 803 31040 890
rect 31040 803 31127 890
rect 31127 803 31133 890
rect 31034 797 31133 803
rect 18113 406 18165 415
rect 18113 372 18122 406
rect 18122 372 18156 406
rect 18156 372 18165 406
rect 18113 363 18165 372
rect 22518 307 22570 316
rect 22518 273 22527 307
rect 22527 273 22561 307
rect 22561 273 22570 307
rect 22518 264 22570 273
rect 26927 306 26979 315
rect 26927 272 26936 306
rect 26936 272 26970 306
rect 26970 272 26979 306
rect 26927 263 26979 272
rect 31347 306 31399 315
rect 31347 272 31356 306
rect 31356 272 31390 306
rect 31390 272 31399 306
rect 31347 263 31399 272
<< metal2 >>
rect 19961 11345 20278 11355
rect 19961 11048 19972 11345
rect 20269 11048 20278 11345
rect 19961 11038 20278 11048
rect 20634 8774 20765 8780
rect 20634 8655 20640 8774
rect 20759 8655 20765 8774
rect 20634 8649 20765 8655
rect 21544 8678 21611 8686
rect 19962 6530 20279 6542
rect 19962 6233 19972 6530
rect 20269 6233 20279 6530
rect 19962 6223 20279 6233
rect 20646 5204 20753 8649
rect 21544 8626 21551 8678
rect 21603 8626 21611 8678
rect 21544 5460 21611 8626
rect 21718 8669 21783 8676
rect 21718 8617 21724 8669
rect 21776 8617 21783 8669
rect 21718 6065 21783 8617
rect 25018 7556 25140 7586
rect 25018 7494 25048 7556
rect 25110 7494 25140 7556
rect 21718 5994 23508 6065
rect 21544 5404 22944 5460
rect 20646 5149 22409 5204
rect 22606 5202 22658 5208
rect 22374 2018 22408 5149
rect 22606 5144 22658 5150
rect 22359 2012 22423 2018
rect 22615 2016 22649 5144
rect 22888 4870 22944 5404
rect 22882 4814 22888 4870
rect 22944 4814 22950 4870
rect 23459 4374 23508 5994
rect 25018 5967 25140 7494
rect 25493 7437 25574 7447
rect 25493 7375 25502 7437
rect 25564 7375 25574 7437
rect 25045 5202 25110 5967
rect 25045 5150 25051 5202
rect 25103 5150 25110 5202
rect 25045 5144 25110 5150
rect 25493 5051 25574 7375
rect 27071 6018 27252 6025
rect 27071 5850 27077 6018
rect 27245 6012 27252 6018
rect 27245 5856 31524 6012
rect 27245 5850 27252 5856
rect 27071 5843 27252 5850
rect 25493 4979 27069 5051
rect 25493 4978 25566 4979
rect 26746 4868 26798 4874
rect 26746 4810 26798 4816
rect 23459 4322 23465 4374
rect 23517 4322 23523 4374
rect 22359 1960 22365 2012
rect 22417 1960 22423 2012
rect 22359 1954 22423 1960
rect 22600 2010 22664 2016
rect 22600 1958 22606 2010
rect 22658 1958 22664 2010
rect 26755 1999 26789 4810
rect 27013 2001 27069 4979
rect 31143 4322 31149 4374
rect 31201 4322 31207 4374
rect 31158 2068 31192 4322
rect 31149 2062 31201 2068
rect 31149 2004 31201 2010
rect 22600 1952 22664 1958
rect 26740 1993 26804 1999
rect 26740 1941 26746 1993
rect 26798 1941 26804 1993
rect 26740 1935 26804 1941
rect 27009 1995 27073 2001
rect 27009 1943 27015 1995
rect 27067 1943 27073 1995
rect 27009 1937 27073 1943
rect 31368 1883 31524 5856
rect 31368 1721 31524 1727
rect 22712 1262 22843 1272
rect 18271 1183 18396 1192
rect 17453 1143 17686 1153
rect 17453 932 17462 1143
rect 17673 932 17686 1143
rect 18271 1071 18277 1183
rect 18389 1071 18396 1183
rect 22712 1149 22721 1262
rect 22834 1149 22843 1262
rect 27120 1270 27250 1279
rect 27120 1158 27129 1270
rect 27241 1158 27250 1270
rect 27120 1149 27250 1158
rect 30849 1255 30979 1264
rect 22712 1140 22843 1149
rect 30849 1143 30858 1255
rect 30970 1143 30979 1255
rect 30849 1134 30979 1143
rect 18271 1065 18396 1071
rect 27294 973 27414 984
rect 17453 923 17686 932
rect 22888 930 23004 941
rect 18444 876 18560 887
rect 16949 800 17161 807
rect 16949 601 16955 800
rect 17154 601 17161 800
rect 18444 778 18453 876
rect 18551 778 18560 876
rect 22888 832 22897 930
rect 22995 832 23004 930
rect 27294 875 27305 973
rect 27403 875 27414 973
rect 27294 864 27414 875
rect 31022 896 31144 907
rect 22888 823 23004 832
rect 31022 797 31034 896
rect 31133 797 31144 896
rect 31022 786 31144 797
rect 18444 768 18560 778
rect 16949 595 17161 601
rect 18086 419 18194 440
rect 18086 359 18109 419
rect 18169 359 18194 419
rect 18086 336 18194 359
rect 22492 320 22594 340
rect 22492 260 22514 320
rect 22574 260 22594 320
rect 22492 244 22594 260
rect 26901 319 27003 339
rect 26901 259 26923 319
rect 26983 259 27003 319
rect 26901 243 27003 259
rect 31321 319 31423 339
rect 31321 259 31343 319
rect 31403 259 31423 319
rect 31321 243 31423 259
<< via2 >>
rect 19972 11048 20269 11345
rect 19972 6233 20269 6530
rect 17462 932 17673 1143
rect 18277 1083 18389 1183
rect 22721 1149 22834 1262
rect 27129 1158 27241 1270
rect 30858 1143 30970 1255
rect 16960 606 17149 795
rect 18453 778 18551 876
rect 22897 832 22995 930
rect 27305 875 27403 973
rect 31034 797 31133 896
rect 18109 415 18169 419
rect 18109 363 18113 415
rect 18113 363 18165 415
rect 18165 363 18169 415
rect 18109 359 18169 363
rect 22514 316 22574 320
rect 22514 264 22518 316
rect 22518 264 22570 316
rect 22570 264 22574 316
rect 22514 260 22574 264
rect 26923 315 26983 319
rect 26923 263 26927 315
rect 26927 263 26979 315
rect 26979 263 26983 315
rect 26923 259 26983 263
rect 31343 315 31403 319
rect 31343 263 31347 315
rect 31347 263 31399 315
rect 31399 263 31403 315
rect 31343 259 31403 263
<< metal3 >>
rect 9794 26731 9800 27131
rect 10200 27130 20105 27131
rect 10200 26732 19706 27130
rect 20104 26732 20110 27130
rect 10200 26731 20105 26732
rect 19967 11345 20274 11350
rect 9801 11048 9807 11345
rect 10104 11048 19972 11345
rect 20269 11048 20274 11345
rect 19967 11043 20274 11048
rect 4224 9101 9919 9229
rect 10047 9101 10053 9229
rect 19967 6530 20274 6535
rect 9794 6233 9800 6530
rect 10097 6233 19972 6530
rect 20269 6233 20274 6530
rect 19967 6228 20274 6233
rect 4057 3742 8732 3743
rect 4057 3564 8553 3742
rect 8731 3564 8737 3742
rect 4057 3563 8732 3564
rect 200 1864 31128 1870
rect 200 1652 243 1864
rect 455 1652 31128 1864
rect 200 1646 31128 1652
rect 9800 1446 16941 1471
rect 9800 1288 9860 1446
rect 10005 1288 16941 1446
rect 9800 1272 16941 1288
rect 17142 1272 17154 1471
rect 16955 795 17154 1272
rect 17462 1148 17686 1646
rect 18283 1192 18383 1646
rect 22727 1267 22828 1646
rect 27135 1275 27235 1646
rect 27124 1270 27246 1275
rect 22716 1262 22839 1267
rect 17457 1143 17686 1148
rect 17457 932 17462 1143
rect 17673 938 17686 1143
rect 18271 1183 18396 1192
rect 18271 1083 18277 1183
rect 18389 1083 18396 1183
rect 22716 1149 22721 1262
rect 22834 1149 22839 1262
rect 27124 1158 27129 1270
rect 27241 1158 27246 1270
rect 30864 1260 30964 1646
rect 27124 1153 27246 1158
rect 30853 1255 30975 1260
rect 22716 1144 22839 1149
rect 30853 1143 30858 1255
rect 30970 1143 30975 1255
rect 30853 1138 30975 1143
rect 18271 1065 18396 1083
rect 27294 978 27414 984
rect 17673 932 17678 938
rect 17457 927 17678 932
rect 22892 935 23000 941
rect 16955 606 16960 795
rect 17149 606 17154 795
rect 18444 881 18560 887
rect 18444 795 18448 881
rect 18556 795 18560 881
rect 27294 870 27300 978
rect 27408 870 27414 978
rect 27294 864 27414 870
rect 31022 901 31144 907
rect 22892 832 22897 849
rect 22995 832 23000 849
rect 22892 827 23000 832
rect 18444 778 18453 795
rect 18551 778 18560 795
rect 31022 792 31029 901
rect 31138 792 31144 901
rect 31022 786 31144 792
rect 18444 768 18560 778
rect 16955 601 17154 606
rect 18086 424 18194 440
rect 18086 354 18104 424
rect 18174 354 18194 424
rect 18086 336 18194 354
rect 22492 325 22594 340
rect 22492 255 22509 325
rect 22579 255 22594 325
rect 22492 244 22594 255
rect 26901 324 27003 339
rect 26901 254 26918 324
rect 26988 254 27003 324
rect 26901 243 27003 254
rect 31321 324 31423 339
rect 31321 254 31338 324
rect 31408 254 31423 324
rect 31321 243 31423 254
<< via3 >>
rect 9800 26731 10200 27131
rect 19706 26732 20104 27130
rect 9807 11048 10104 11345
rect 9919 9101 10047 9229
rect 9800 6233 10097 6530
rect 8553 3564 8731 3742
rect 243 1652 455 1864
rect 9860 1288 10005 1446
rect 16941 1272 17142 1471
rect 22892 930 23000 935
rect 18448 876 18556 881
rect 18448 795 18453 876
rect 18453 795 18551 876
rect 18551 795 18556 876
rect 22892 849 22897 930
rect 22897 849 22995 930
rect 22995 849 23000 930
rect 27300 973 27408 978
rect 27300 875 27305 973
rect 27305 875 27403 973
rect 27403 875 27408 973
rect 27300 870 27408 875
rect 31029 896 31138 901
rect 31029 797 31034 896
rect 31034 797 31133 896
rect 31133 797 31138 896
rect 31029 792 31138 797
rect 18104 419 18174 424
rect 18104 359 18109 419
rect 18109 359 18169 419
rect 18169 359 18174 419
rect 18104 354 18174 359
rect 22509 320 22579 325
rect 22509 260 22514 320
rect 22514 260 22574 320
rect 22574 260 22579 320
rect 22509 255 22579 260
rect 26918 319 26988 324
rect 26918 259 26923 319
rect 26923 259 26983 319
rect 26983 259 26988 319
rect 26918 254 26988 259
rect 31338 319 31408 324
rect 31338 259 31343 319
rect 31343 259 31403 319
rect 31403 259 31408 319
rect 31338 254 31408 259
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 1864 500 44152
rect 9800 27132 10100 44152
rect 9799 27131 10201 27132
rect 9799 26731 9800 27131
rect 10200 26731 10201 27131
rect 9799 26730 10201 26731
rect 9800 11346 10100 26730
rect 18905 25955 19305 28937
rect 19705 27130 20105 28565
rect 19705 26732 19706 27130
rect 20104 26732 20105 27130
rect 19705 26731 20105 26732
rect 11538 25555 19305 25955
rect 9800 11345 10105 11346
rect 9800 11048 9807 11345
rect 10104 11048 10105 11345
rect 9800 11047 10105 11048
rect 9800 9229 10100 11047
rect 9800 9101 9919 9229
rect 10047 9101 10100 9229
rect 9800 6531 10100 9101
rect 9799 6530 10100 6531
rect 9799 6233 9800 6530
rect 10097 6233 10100 6530
rect 9799 6232 10100 6233
rect 200 1652 243 1864
rect 455 1652 500 1864
rect 200 1000 500 1652
rect 8552 3742 8732 3743
rect 8552 3564 8553 3742
rect 8731 3564 8732 3742
rect 8552 200 8732 3564
rect 9800 1446 10100 6232
rect 9800 1288 9860 1446
rect 10005 1288 10100 1446
rect 9800 1000 10100 1288
rect 11538 1050 11938 25555
rect 16940 1471 17143 1472
rect 16940 1272 16941 1471
rect 17142 1272 31127 1471
rect 16940 1271 17143 1272
rect 11538 650 13798 1050
rect 18459 887 18545 1272
rect 22903 936 22989 1272
rect 27311 979 27397 1272
rect 27299 978 27409 979
rect 22891 935 23001 936
rect 18444 881 18560 887
rect 18444 795 18448 881
rect 18556 795 18560 881
rect 22891 849 22892 935
rect 23000 849 23001 935
rect 27299 870 27300 978
rect 27408 870 27409 978
rect 31040 902 31127 1272
rect 27299 869 27409 870
rect 31028 901 31139 902
rect 22891 848 23001 849
rect 18444 768 18560 795
rect 31028 792 31029 901
rect 31138 792 31139 901
rect 31028 791 31139 792
rect 370 0 550 200
rect 4786 0 4966 200
rect 8552 20 9382 200
rect 9202 0 9382 20
rect 13618 0 13798 650
rect 18086 424 18194 440
rect 18086 354 18104 424
rect 18174 354 18194 424
rect 18086 336 18194 354
rect 18109 200 18169 336
rect 22492 325 22594 340
rect 22492 255 22509 325
rect 22579 255 22594 325
rect 22492 200 22594 255
rect 26901 324 27003 339
rect 26901 254 26918 324
rect 26988 254 27003 324
rect 26901 200 27003 254
rect 31321 324 31423 339
rect 31321 254 31338 324
rect 31408 254 31423 324
rect 31321 200 31423 254
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use bodynmos  bodynmos_0
timestamp 1716541817
transform 1 0 22927 0 1 777
box -24 -24 62 52
use bodynmos  bodynmos_1
timestamp 1716541817
transform 1 0 18483 0 1 688
box -24 -24 62 52
use bodynmos  bodynmos_2
timestamp 1716541817
transform 1 0 27335 0 1 775
box -24 -24 62 52
use bodynmos  bodynmos_3
timestamp 1716541817
transform 1 0 31064 0 1 738
box -24 -24 62 52
use bodypmos  bodypmos_0
timestamp 1716540843
transform 1 0 22765 0 1 1111
box -76 -78 118 110
use bodypmos  bodypmos_1
timestamp 1716540843
transform 1 0 18321 0 1 1022
box -76 -78 118 110
use bodypmos  bodypmos_2
timestamp 1716540843
transform 1 0 27173 0 1 1109
box -76 -78 118 110
use bodypmos  bodypmos_3
timestamp 1716540843
transform 1 0 30902 0 1 1056
box -76 -78 118 110
use compschematic  compschematic_0
timestamp 1717263723
transform 1 0 21047 0 1 8570
box -314 -358 510 960
use inductor  inductor_0
timestamp 1717235020
transform 1 0 3844 0 1 3873
box 0 -412 510 5490
use inverter  inverter_0
timestamp 1717263723
transform 1 0 18078 0 1 -67
box -226 644 170 1266
use loop_antenna  loop_antenna_0
timestamp 1717233969
transform 1 0 19705 0 -1 34537
box -5000 -8800 8200 6000
use mux1_2  mux1_2_0
timestamp 1717263723
transform 1 0 31220 0 1 527
box 0 98 306 776
use mux1_2  mux1_2_3
timestamp 1717263723
transform 1 0 22391 0 1 528
box 0 98 306 776
use mux1_2  mux1_2_4
timestamp 1717263723
transform 1 0 26800 0 1 527
box 0 98 306 776
use new_latest  new_latest_0
timestamp 1717250560
transform 1 0 27281 0 1 5875
box -3192 359 1303 5470
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
