magic
tech sky130A
magscale 1 2
timestamp 1716458959
<< metal3 >>
rect -386 3092 386 3120
rect -386 2668 302 3092
rect 366 2668 386 3092
rect -386 2640 386 2668
rect -386 2372 386 2400
rect -386 1948 302 2372
rect 366 1948 386 2372
rect -386 1920 386 1948
rect -386 1652 386 1680
rect -386 1228 302 1652
rect 366 1228 386 1652
rect -386 1200 386 1228
rect -386 932 386 960
rect -386 508 302 932
rect 366 508 386 932
rect -386 480 386 508
rect -386 212 386 240
rect -386 -212 302 212
rect 366 -212 386 212
rect -386 -240 386 -212
rect -386 -508 386 -480
rect -386 -932 302 -508
rect 366 -932 386 -508
rect -386 -960 386 -932
rect -386 -1228 386 -1200
rect -386 -1652 302 -1228
rect 366 -1652 386 -1228
rect -386 -1680 386 -1652
rect -386 -1948 386 -1920
rect -386 -2372 302 -1948
rect 366 -2372 386 -1948
rect -386 -2400 386 -2372
rect -386 -2668 386 -2640
rect -386 -3092 302 -2668
rect 366 -3092 386 -2668
rect -386 -3120 386 -3092
<< via3 >>
rect 302 2668 366 3092
rect 302 1948 366 2372
rect 302 1228 366 1652
rect 302 508 366 932
rect 302 -212 366 212
rect 302 -932 366 -508
rect 302 -1652 366 -1228
rect 302 -2372 366 -1948
rect 302 -3092 366 -2668
<< mimcap >>
rect -346 3040 54 3080
rect -346 2720 -306 3040
rect 14 2720 54 3040
rect -346 2680 54 2720
rect -346 2320 54 2360
rect -346 2000 -306 2320
rect 14 2000 54 2320
rect -346 1960 54 2000
rect -346 1600 54 1640
rect -346 1280 -306 1600
rect 14 1280 54 1600
rect -346 1240 54 1280
rect -346 880 54 920
rect -346 560 -306 880
rect 14 560 54 880
rect -346 520 54 560
rect -346 160 54 200
rect -346 -160 -306 160
rect 14 -160 54 160
rect -346 -200 54 -160
rect -346 -560 54 -520
rect -346 -880 -306 -560
rect 14 -880 54 -560
rect -346 -920 54 -880
rect -346 -1280 54 -1240
rect -346 -1600 -306 -1280
rect 14 -1600 54 -1280
rect -346 -1640 54 -1600
rect -346 -2000 54 -1960
rect -346 -2320 -306 -2000
rect 14 -2320 54 -2000
rect -346 -2360 54 -2320
rect -346 -2720 54 -2680
rect -346 -3040 -306 -2720
rect 14 -3040 54 -2720
rect -346 -3080 54 -3040
<< mimcapcontact >>
rect -306 2720 14 3040
rect -306 2000 14 2320
rect -306 1280 14 1600
rect -306 560 14 880
rect -306 -160 14 160
rect -306 -880 14 -560
rect -306 -1600 14 -1280
rect -306 -2320 14 -2000
rect -306 -3040 14 -2720
<< metal4 >>
rect -198 3041 -94 3240
rect 282 3092 386 3240
rect -307 3040 15 3041
rect -307 2720 -306 3040
rect 14 2720 15 3040
rect -307 2719 15 2720
rect -198 2321 -94 2719
rect 282 2668 302 3092
rect 366 2668 386 3092
rect 282 2372 386 2668
rect -307 2320 15 2321
rect -307 2000 -306 2320
rect 14 2000 15 2320
rect -307 1999 15 2000
rect -198 1601 -94 1999
rect 282 1948 302 2372
rect 366 1948 386 2372
rect 282 1652 386 1948
rect -307 1600 15 1601
rect -307 1280 -306 1600
rect 14 1280 15 1600
rect -307 1279 15 1280
rect -198 881 -94 1279
rect 282 1228 302 1652
rect 366 1228 386 1652
rect 282 932 386 1228
rect -307 880 15 881
rect -307 560 -306 880
rect 14 560 15 880
rect -307 559 15 560
rect -198 161 -94 559
rect 282 508 302 932
rect 366 508 386 932
rect 282 212 386 508
rect -307 160 15 161
rect -307 -160 -306 160
rect 14 -160 15 160
rect -307 -161 15 -160
rect -198 -559 -94 -161
rect 282 -212 302 212
rect 366 -212 386 212
rect 282 -508 386 -212
rect -307 -560 15 -559
rect -307 -880 -306 -560
rect 14 -880 15 -560
rect -307 -881 15 -880
rect -198 -1279 -94 -881
rect 282 -932 302 -508
rect 366 -932 386 -508
rect 282 -1228 386 -932
rect -307 -1280 15 -1279
rect -307 -1600 -306 -1280
rect 14 -1600 15 -1280
rect -307 -1601 15 -1600
rect -198 -1999 -94 -1601
rect 282 -1652 302 -1228
rect 366 -1652 386 -1228
rect 282 -1948 386 -1652
rect -307 -2000 15 -1999
rect -307 -2320 -306 -2000
rect 14 -2320 15 -2000
rect -307 -2321 15 -2320
rect -198 -2719 -94 -2321
rect 282 -2372 302 -1948
rect 366 -2372 386 -1948
rect 282 -2668 386 -2372
rect -307 -2720 15 -2719
rect -307 -3040 -306 -2720
rect 14 -3040 15 -2720
rect -307 -3041 15 -3040
rect -198 -3240 -94 -3041
rect 282 -3092 302 -2668
rect 366 -3092 386 -2668
rect 282 -3240 386 -3092
<< properties >>
string FIXED_BBOX -386 2640 94 3120
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 9 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
