magic
tech sky130A
timestamp 1717240620
<< pwell >>
rect -198 -455 198 455
<< nmos >>
rect -100 -350 100 350
<< ndiff >>
rect -129 344 -100 350
rect -129 -344 -123 344
rect -106 -344 -100 344
rect -129 -350 -100 -344
rect 100 344 129 350
rect 100 -344 106 344
rect 123 -344 129 344
rect 100 -350 129 -344
<< ndiffc >>
rect -123 -344 -106 344
rect 106 -344 123 344
<< psubdiff >>
rect -180 420 -132 437
rect 132 420 180 437
rect -180 389 -163 420
rect 163 389 180 420
rect -180 -420 -163 -389
rect 163 -420 180 -389
rect -180 -437 -132 -420
rect 132 -437 180 -420
<< psubdiffcont >>
rect -132 420 132 437
rect -180 -389 -163 389
rect 163 -389 180 389
rect -132 -437 132 -420
<< poly >>
rect -100 386 100 394
rect -100 369 -92 386
rect 92 369 100 386
rect -100 350 100 369
rect -100 -369 100 -350
rect -100 -386 -92 -369
rect 92 -386 100 -369
rect -100 -394 100 -386
<< polycont >>
rect -92 369 92 386
rect -92 -386 92 -369
<< locali >>
rect -180 420 -132 437
rect 132 420 180 437
rect -180 389 -163 420
rect 163 389 180 420
rect -100 369 -92 386
rect 92 369 100 386
rect -123 344 -106 352
rect -123 -352 -106 -344
rect 106 344 123 352
rect 106 -352 123 -344
rect -100 -386 -92 -369
rect 92 -386 100 -369
rect -180 -420 -163 -389
rect 163 -420 180 -389
rect -180 -437 -132 -420
rect 132 -437 180 -420
<< viali >>
rect -92 369 92 386
rect -123 -344 -106 344
rect 106 -344 123 344
rect -92 -386 92 -369
<< metal1 >>
rect -98 386 98 389
rect -98 369 -92 386
rect 92 369 98 386
rect -98 366 98 369
rect -126 344 -103 350
rect -126 -344 -123 344
rect -106 -344 -103 344
rect -126 -350 -103 -344
rect 103 344 126 350
rect 103 -344 106 344
rect 123 -344 126 344
rect 103 -350 126 -344
rect -98 -369 98 -366
rect -98 -386 -92 -369
rect 92 -386 98 -369
rect -98 -389 98 -386
<< properties >>
string FIXED_BBOX -171 -428 171 428
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 7.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
